-------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
-------------------------------------------------------------------------------
-- Generated from "TEST80.BIN"
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Package with utility functions for handling SoC object code.
use work.mcu80_pkg.all;

package obj_code_pkg is

-- Object code initialization constant.
constant object_code : obj_code_t(0 to 16383) := (
  X"31",X"00",X"00",X"3e",X"00",X"32",X"00",X"f8", -- 0000
  X"32",X"01",X"f8",X"32",X"02",X"f8",X"d3",X"01", -- 0008
  X"d3",X"01",X"d3",X"01",X"3e",X"40",X"d3",X"01", -- 0010
  X"3e",X"4e",X"d3",X"01",X"3e",X"37",X"d3",X"01", -- 0018
  X"fb",X"c3",X"8d",X"00",X"f5",X"db",X"01",X"e6", -- 0020
  X"01",X"ca",X"25",X"00",X"f1",X"d3",X"00",X"c9", -- 0028
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0030
  X"f3",X"f5",X"c5",X"d5",X"e5",X"db",X"01",X"e6", -- 0038
  X"02",X"ca",X"62",X"00",X"db",X"00",X"57",X"3a", -- 0040
  X"00",X"f8",X"fe",X"ff",X"ca",X"62",X"00",X"3c", -- 0048
  X"32",X"00",X"f8",X"3a",X"02",X"f8",X"4f",X"06", -- 0050
  X"00",X"21",X"03",X"f8",X"09",X"72",X"3c",X"32", -- 0058
  X"02",X"f8",X"e1",X"d1",X"c1",X"f1",X"fb",X"c9", -- 0060
  X"c5",X"d5",X"e5",X"3a",X"00",X"f8",X"fe",X"00", -- 0068
  X"ca",X"6b",X"00",X"f3",X"3d",X"32",X"00",X"f8", -- 0070
  X"3a",X"01",X"f8",X"4f",X"06",X"00",X"21",X"03", -- 0078
  X"f8",X"09",X"56",X"3c",X"32",X"01",X"f8",X"7a", -- 0080
  X"fb",X"e1",X"d1",X"c1",X"c9",X"3e",X"3e",X"cd", -- 0088
  X"24",X"00",X"cd",X"68",X"00",X"cd",X"24",X"00", -- 0090
  X"c3",X"92",X"00",X"00",X"00",X"00",X"00",X"00", -- 0098
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 00f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0100
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0108
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0110
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0118
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0120
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0128
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0130
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0138
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0140
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0148
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0150
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0158
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0160
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0168
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0170
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0178
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0180
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0188
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0190
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0198
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 01f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0200
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0208
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0210
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0218
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0220
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0228
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0230
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0238
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0240
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0248
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0250
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0258
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0260
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0268
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0270
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0278
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0280
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0288
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0290
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0298
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 02f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0300
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0308
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0310
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0318
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0320
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0328
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0330
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0338
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0340
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0348
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0350
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0358
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0360
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0368
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0370
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0378
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0380
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0388
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0390
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0398
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 03f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0400
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0408
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0410
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0418
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0420
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0428
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0430
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0438
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0440
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0448
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0450
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0458
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0460
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0468
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0470
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0478
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0480
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0488
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0490
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0498
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 04f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0500
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0508
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0510
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0518
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0520
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0528
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0530
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0538
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0540
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0548
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0550
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0558
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0560
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0568
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0570
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0578
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0580
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0588
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0590
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0598
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 05f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0600
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0608
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0610
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0618
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0620
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0628
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0630
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0638
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0640
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0648
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0650
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0658
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0660
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0668
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0670
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0678
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0680
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0688
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0690
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0698
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 06f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0700
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0708
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0710
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0718
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0720
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0728
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0730
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0738
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0740
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0748
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0750
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0758
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0760
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0768
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0770
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0778
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0780
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0788
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0790
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0798
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 07f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0800
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0808
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0810
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0818
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0820
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0828
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0830
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0838
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0840
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0848
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0850
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0858
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0860
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0868
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0870
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0878
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0880
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0888
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0890
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0898
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 08f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0900
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0908
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0910
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0918
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0920
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0928
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0930
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0938
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0940
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0948
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0950
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0958
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0960
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0968
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0970
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0978
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0980
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0988
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0990
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0998
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 09f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0a98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0aa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0aa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ab0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ab8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ac0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ac8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ad0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ad8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ae0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ae8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0af0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0af8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0b98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ba0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ba8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0bb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0bb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0bc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0bc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0bd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0bd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0be0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0be8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0bf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0bf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0c98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ca0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ca8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0cb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0cb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0cc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0cc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0cd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0cd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ce0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ce8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0cf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0cf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0d98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0da0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0da8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0db0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0db8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0dc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0dc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0dd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0dd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0de0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0de8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0df0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0df8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0e98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ea0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ea8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0eb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0eb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ec0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ec8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ed0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ed8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ee0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ee8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ef0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ef8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0f98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0fa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0fa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0fb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0fb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0fc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0fc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0fd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0fd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0fe0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0fe8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ff0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0ff8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1000
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1008
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1010
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1018
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1020
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1028
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1030
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1038
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1040
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1048
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1050
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1058
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1060
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1068
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1070
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1078
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1080
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1088
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1090
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1098
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1100
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1108
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1110
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1118
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1120
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1128
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1130
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1138
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1140
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1148
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1150
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1158
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1160
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1168
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1170
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1178
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1180
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1188
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1190
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1198
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1200
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1208
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1210
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1218
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1220
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1228
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1230
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1238
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1240
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1248
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1250
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1258
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1260
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1268
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1270
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1278
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1280
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1288
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1290
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1298
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1300
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1308
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1310
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1318
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1320
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1328
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1330
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1338
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1340
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1348
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1350
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1358
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1360
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1368
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1370
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1378
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1380
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1388
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1390
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1398
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1400
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1408
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1410
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1418
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1420
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1428
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1430
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1438
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1440
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1448
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1450
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1458
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1460
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1468
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1470
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1478
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1480
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1488
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1490
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1498
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 14f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1500
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1508
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1510
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1518
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1520
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1528
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1530
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1538
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1540
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1548
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1550
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1558
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1560
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1568
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1570
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1578
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1580
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1588
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1590
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1598
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 15f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1600
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1608
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1610
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1618
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1620
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1628
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1630
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1638
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1640
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1648
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1650
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1658
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1660
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1668
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1670
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1678
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1680
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1688
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1690
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1698
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 16f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1700
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1708
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1710
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1718
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1720
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1728
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1730
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1738
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1740
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1748
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1750
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1758
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1760
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1768
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1770
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1778
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1780
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1788
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1790
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1798
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 17f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1800
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1808
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1810
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1818
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1820
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1828
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1830
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1838
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1840
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1848
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1850
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1858
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1860
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1868
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1870
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1878
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1880
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1888
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1890
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1898
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 18f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1900
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1908
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1910
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1918
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1920
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1928
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1930
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1938
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1940
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1948
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1950
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1958
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1960
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1968
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1970
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1978
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1980
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1988
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1990
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1998
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 19f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1a98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1aa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1aa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ab0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ab8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ac0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ac8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ad0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ad8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ae0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ae8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1af0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1af8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1b98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ba0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ba8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1bb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1bb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1bc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1bc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1bd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1bd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1be0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1be8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1bf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1bf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1c98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ca0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ca8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1cb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1cb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1cc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1cc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1cd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1cd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ce0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ce8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1cf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1cf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1da0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1da8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1db0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1db8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1dc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1dc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1dd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1dd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1de0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1de8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1df0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1df8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ea0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ea8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1eb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1eb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ec0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ec8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ed0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ed8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ee0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ee8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ef0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ef8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fe0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fe8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ff0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ff8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2000
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2008
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2010
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2018
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2020
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2028
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2030
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2038
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2040
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2048
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2050
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2058
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2060
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2068
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2070
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2078
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2080
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2088
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2090
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2098
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2100
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2108
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2110
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2118
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2120
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2128
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2130
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2138
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2140
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2148
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2150
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2158
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2160
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2168
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2170
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2178
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2180
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2188
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2190
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2198
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2200
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2208
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2210
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2218
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2220
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2228
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2230
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2238
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2240
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2248
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2250
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2258
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2260
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2268
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2270
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2278
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2280
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2288
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2290
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2298
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2300
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2308
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2310
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2318
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2320
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2328
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2330
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2338
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2340
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2348
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2350
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2358
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2360
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2368
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2370
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2378
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2380
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2388
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2390
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2398
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2400
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2408
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2410
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2418
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2420
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2428
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2430
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2438
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2440
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2448
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2450
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2458
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2460
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2468
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2470
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2478
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2480
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2488
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2490
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2498
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2500
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2508
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2510
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2518
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2520
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2528
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2530
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2538
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2540
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2548
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2550
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2558
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2560
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2568
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2570
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2578
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2580
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2588
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2590
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2598
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2600
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2608
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2610
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2618
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2620
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2628
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2630
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2638
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2640
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2648
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2650
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2658
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2660
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2668
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2670
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2678
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2680
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2688
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2690
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2698
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2700
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2708
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2710
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2718
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2720
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2728
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2730
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2738
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2740
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2748
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2750
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2758
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2760
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2768
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2770
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2778
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2780
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2788
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2790
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2798
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2800
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2808
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2810
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2818
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2820
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2828
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2830
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2838
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2840
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2848
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2850
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2858
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2860
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2868
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2870
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2878
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2880
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2888
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2890
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2898
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2900
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2908
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2910
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2918
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2920
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2928
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2930
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2938
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2940
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2948
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2950
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2958
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2960
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2968
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2970
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2978
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2980
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2988
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2990
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2998
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2aa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2aa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ab0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ab8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ac0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ac8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ad0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ad8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ae0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ae8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2af0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2af8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ba0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ba8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2be0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2be8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ca0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ca8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ce0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ce8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2da0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2da8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2db0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2db8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2de0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2de8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2df0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2df8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ea0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ea8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2eb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2eb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ec0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ec8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ed0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ed8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ee0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ee8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ef0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ef8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fe0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fe8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ff0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ff8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3000
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3008
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3010
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3018
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3020
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3028
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3030
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3038
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3040
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3048
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3050
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3058
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3060
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3068
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3070
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3078
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3080
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3088
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3090
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3098
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3100
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3108
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3110
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3118
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3120
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3128
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3130
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3138
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3140
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3148
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3150
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3158
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3160
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3168
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3170
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3178
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3180
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3188
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3190
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3198
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3200
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3208
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3210
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3218
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3220
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3228
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3230
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3238
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3240
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3248
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3250
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3258
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3260
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3268
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3270
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3278
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3280
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3288
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3290
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3298
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3300
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3308
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3310
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3318
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3320
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3328
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3330
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3338
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3340
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3348
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3350
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3358
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3360
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3368
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3370
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3378
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3380
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3388
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3390
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3398
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3400
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3408
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3410
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3418
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3420
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3428
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3430
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3438
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3440
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3448
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3450
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3458
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3460
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3468
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3470
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3478
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3480
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3488
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3490
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3498
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3500
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3508
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3510
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3518
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3520
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3528
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3530
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3538
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3540
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3548
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3550
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3558
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3560
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3568
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3570
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3578
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3580
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3588
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3590
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3598
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3600
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3608
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3610
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3618
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3620
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3628
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3630
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3638
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3640
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3648
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3650
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3658
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3660
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3668
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3670
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3678
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3680
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3688
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3690
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3698
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3700
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3708
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3710
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3718
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3720
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3728
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3730
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3738
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3740
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3748
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3750
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3758
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3760
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3768
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3770
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3778
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3780
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3788
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3790
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3798
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3800
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3808
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3810
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3818
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3820
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3828
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3830
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3838
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3840
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3848
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3850
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3858
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3860
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3868
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3870
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3878
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3880
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3888
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3890
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3898
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3900
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3908
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3910
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3918
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3920
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3928
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3930
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3938
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3940
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3948
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3950
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3958
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3960
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3968
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3970
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3978
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3980
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3988
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3990
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3998
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3aa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3aa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ab0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ab8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ac0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ac8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ad0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ad8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ae0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ae8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3af0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3af8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ba0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ba8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3be0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3be8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ca0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ca8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ce0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ce8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3da0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3da8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3db0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3db8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3de0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3de8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3df0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3df8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ea0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ea8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3eb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3eb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ec0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ec8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ed0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ed8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ee0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ee8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ef0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ef8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fe0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fe8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ff0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"  -- 3ff8
  );

end package obj_code_pkg;
