-------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
-------------------------------------------------------------------------------
-- Generated from "MON80SA.BIN"
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Package with utility functions for handling SoC object code.
use work.mcu80_pkg.all;

package obj_code_pkg is

-- Object code initialization constant.
constant object_code : obj_code_t(0 to 16383) := (
  X"c3",X"d4",X"00",X"00",X"00",X"f5",X"79",X"07", -- 0000
  X"81",X"4f",X"f1",X"06",X"00",X"21",X"12",X"00", -- 0008
  X"09",X"e9",X"c3",X"d4",X"00",X"c3",X"7c",X"00", -- 0010
  X"c3",X"ab",X"00",X"c3",X"7c",X"00",X"c3",X"ab", -- 0018
  X"00",X"c3",X"ab",X"00",X"c3",X"c0",X"00",X"db", -- 0020
  X"01",X"e6",X"02",X"ca",X"27",X"00",X"db",X"00", -- 0028
  X"c9",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0030
  X"f3",X"f5",X"c5",X"d5",X"e5",X"cd",X"27",X"00", -- 0038
  X"fe",X"11",X"ca",X"4a",X"00",X"fe",X"13",X"c2", -- 0040
  X"50",X"00",X"32",X"ff",X"fe",X"c3",X"76",X"00", -- 0048
  X"57",X"3a",X"fc",X"fe",X"fe",X"ff",X"ca",X"76", -- 0050
  X"00",X"fe",X"af",X"c2",X"63",X"00",X"1e",X"13", -- 0058
  X"cd",X"ab",X"00",X"3c",X"32",X"fc",X"fe",X"3a", -- 0060
  X"fe",X"fe",X"4f",X"06",X"00",X"21",X"00",X"ff", -- 0068
  X"09",X"72",X"3c",X"32",X"fe",X"fe",X"e1",X"d1", -- 0070
  X"c1",X"f1",X"fb",X"c9",X"c5",X"d5",X"e5",X"3a", -- 0078
  X"fc",X"fe",X"fe",X"00",X"ca",X"7f",X"00",X"f3", -- 0080
  X"fe",X"af",X"c2",X"92",X"00",X"1e",X"11",X"cd", -- 0088
  X"ab",X"00",X"3d",X"32",X"fc",X"fe",X"3a",X"fd", -- 0090
  X"fe",X"4f",X"06",X"00",X"21",X"00",X"ff",X"09", -- 0098
  X"56",X"3c",X"32",X"fd",X"fe",X"7a",X"fb",X"e1", -- 00a0
  X"d1",X"c1",X"c9",X"f5",X"3a",X"ff",X"fe",X"fe", -- 00a8
  X"13",X"ca",X"ac",X"00",X"db",X"01",X"e6",X"01", -- 00b0
  X"ca",X"b4",X"00",X"7b",X"d3",X"00",X"f1",X"c9", -- 00b8
  X"f5",X"7b",X"fe",X"ff",X"ca",X"ca",X"00",X"c3", -- 00c0
  X"b4",X"00",X"f1",X"3a",X"fc",X"fe",X"fe",X"00", -- 00c8
  X"c8",X"c3",X"7c",X"00",X"31",X"fc",X"fe",X"3e", -- 00d0
  X"11",X"32",X"ff",X"fe",X"3e",X"00",X"32",X"fc", -- 00d8
  X"fe",X"32",X"fd",X"fe",X"32",X"fe",X"fe",X"d3", -- 00e0
  X"01",X"d3",X"01",X"d3",X"01",X"3e",X"40",X"d3", -- 00e8
  X"01",X"3e",X"4e",X"d3",X"01",X"3e",X"37",X"d3", -- 00f0
  X"01",X"3e",X"1d",X"fb",X"c3",X"ff",X"00",X"21", -- 00f8
  X"1c",X"fe",X"39",X"f9",X"21",X"e2",X"01",X"39", -- 0100
  X"eb",X"21",X"00",X"80",X"cd",X"15",X"28",X"21", -- 0108
  X"90",X"01",X"39",X"e5",X"21",X"42",X"01",X"39", -- 0110
  X"e5",X"21",X"f4",X"00",X"39",X"e5",X"21",X"a6", -- 0118
  X"00",X"39",X"e5",X"21",X"58",X"00",X"39",X"e5", -- 0120
  X"21",X"0a",X"00",X"39",X"eb",X"21",X"00",X"00", -- 0128
  X"7d",X"12",X"d1",X"7d",X"12",X"d1",X"7d",X"12", -- 0130
  X"d1",X"7d",X"12",X"d1",X"7d",X"12",X"d1",X"7d", -- 0138
  X"12",X"af",X"cd",X"5c",X"1c",X"21",X"3a",X"04", -- 0140
  X"e5",X"3e",X"01",X"cd",X"ef",X"1d",X"c1",X"af", -- 0148
  X"cd",X"5c",X"1c",X"21",X"5c",X"04",X"e5",X"3e", -- 0150
  X"01",X"cd",X"ef",X"1d",X"c1",X"af",X"cd",X"5c", -- 0158
  X"1c",X"21",X"76",X"04",X"e5",X"3e",X"01",X"cd", -- 0160
  X"ef",X"1d",X"c1",X"af",X"cd",X"5c",X"1c",X"af", -- 0168
  X"cd",X"5c",X"1c",X"21",X"e2",X"01",X"39",X"cd", -- 0170
  X"d5",X"27",X"e5",X"3e",X"01",X"cd",X"96",X"11", -- 0178
  X"c1",X"21",X"90",X"01",X"39",X"e5",X"21",X"49", -- 0180
  X"00",X"e5",X"3e",X"02",X"cd",X"17",X"1e",X"c1", -- 0188
  X"c1",X"21",X"90",X"01",X"39",X"e5",X"21",X"42", -- 0190
  X"01",X"39",X"e5",X"21",X"a4",X"00",X"39",X"e5", -- 0198
  X"3e",X"03",X"cd",X"b6",X"11",X"c1",X"c1",X"c1", -- 01a0
  X"21",X"a0",X"00",X"39",X"e5",X"21",X"52",X"00", -- 01a8
  X"39",X"e5",X"21",X"04",X"00",X"39",X"e5",X"3e", -- 01b0
  X"03",X"cd",X"35",X"13",X"c1",X"c1",X"c1",X"21", -- 01b8
  X"90",X"01",X"39",X"cd",X"c8",X"27",X"7c",X"b5", -- 01c0
  X"ca",X"dc",X"01",X"21",X"f0",X"00",X"39",X"e5", -- 01c8
  X"21",X"42",X"01",X"39",X"e5",X"3e",X"02",X"cd", -- 01d0
  X"28",X"17",X"c1",X"c1",X"21",X"f0",X"00",X"39", -- 01d8
  X"e5",X"21",X"90",X"04",X"e5",X"3e",X"02",X"cd", -- 01e0
  X"54",X"17",X"c1",X"c1",X"7c",X"b5",X"c2",X"73", -- 01e8
  X"02",X"21",X"50",X"00",X"39",X"e5",X"3e",X"01", -- 01f0
  X"cd",X"07",X"16",X"c1",X"7c",X"b5",X"ca",X"15", -- 01f8
  X"02",X"21",X"e2",X"01",X"39",X"e5",X"21",X"52", -- 0200
  X"00",X"39",X"e5",X"3e",X"01",X"cd",X"22",X"1b", -- 0208
  X"c1",X"d1",X"cd",X"15",X"28",X"21",X"00",X"00", -- 0210
  X"39",X"e5",X"3e",X"01",X"cd",X"07",X"16",X"c1", -- 0218
  X"7c",X"b5",X"ca",X"3c",X"02",X"21",X"e0",X"01", -- 0220
  X"39",X"e5",X"21",X"02",X"00",X"39",X"e5",X"3e", -- 0228
  X"01",X"cd",X"22",X"1b",X"c1",X"d1",X"cd",X"15", -- 0230
  X"28",X"c3",X"50",X"02",X"21",X"e0",X"01",X"39", -- 0238
  X"e5",X"21",X"e4",X"01",X"39",X"cd",X"d5",X"27", -- 0240
  X"11",X"10",X"00",X"19",X"d1",X"cd",X"15",X"28", -- 0248
  X"21",X"e2",X"01",X"39",X"e5",X"21",X"e4",X"01", -- 0250
  X"39",X"cd",X"d5",X"27",X"e5",X"21",X"e4",X"01", -- 0258
  X"39",X"cd",X"d5",X"27",X"e5",X"3e",X"02",X"cd", -- 0260
  X"b9",X"04",X"c1",X"c1",X"d1",X"cd",X"15",X"28", -- 0268
  X"c3",X"31",X"04",X"21",X"f0",X"00",X"39",X"e5", -- 0270
  X"21",X"95",X"04",X"e5",X"3e",X"02",X"cd",X"54", -- 0278
  X"17",X"c1",X"c1",X"7c",X"b5",X"c2",X"05",X"03", -- 0280
  X"21",X"50",X"00",X"39",X"e5",X"3e",X"01",X"cd", -- 0288
  X"07",X"16",X"c1",X"7c",X"b5",X"ca",X"ac",X"02", -- 0290
  X"21",X"e2",X"01",X"39",X"e5",X"21",X"52",X"00", -- 0298
  X"39",X"e5",X"3e",X"01",X"cd",X"22",X"1b",X"c1", -- 02a0
  X"d1",X"cd",X"15",X"28",X"21",X"00",X"00",X"39", -- 02a8
  X"e5",X"3e",X"01",X"cd",X"07",X"16",X"c1",X"7c", -- 02b0
  X"b5",X"ca",X"d3",X"02",X"21",X"e0",X"01",X"39", -- 02b8
  X"e5",X"21",X"02",X"00",X"39",X"e5",X"3e",X"01", -- 02c0
  X"cd",X"22",X"1b",X"c1",X"d1",X"cd",X"15",X"28", -- 02c8
  X"c3",X"e2",X"02",X"21",X"e0",X"01",X"39",X"eb", -- 02d0
  X"21",X"e2",X"01",X"39",X"cd",X"d5",X"27",X"cd", -- 02d8
  X"15",X"28",X"21",X"e2",X"01",X"39",X"e5",X"21", -- 02e0
  X"e4",X"01",X"39",X"cd",X"d5",X"27",X"e5",X"21", -- 02e8
  X"e4",X"01",X"39",X"cd",X"d5",X"27",X"e5",X"3e", -- 02f0
  X"02",X"cd",X"0a",X"07",X"c1",X"c1",X"d1",X"cd", -- 02f8
  X"15",X"28",X"c3",X"31",X"04",X"21",X"40",X"01", -- 0300
  X"39",X"cd",X"c8",X"27",X"7c",X"b5",X"c2",X"14", -- 0308
  X"03",X"c3",X"31",X"04",X"21",X"40",X"01",X"39", -- 0310
  X"e5",X"21",X"9a",X"04",X"e5",X"3e",X"02",X"cd", -- 0318
  X"54",X"17",X"c1",X"c1",X"7c",X"b5",X"c2",X"30", -- 0320
  X"03",X"af",X"cd",X"64",X"1f",X"c3",X"31",X"04", -- 0328
  X"21",X"40",X"01",X"39",X"e5",X"21",X"a1",X"04", -- 0330
  X"e5",X"3e",X"02",X"cd",X"54",X"17",X"c1",X"c1", -- 0338
  X"7c",X"b5",X"c2",X"53",X"03",X"21",X"a0",X"00", -- 0340
  X"39",X"e5",X"3e",X"01",X"cd",X"05",X"0a",X"c1", -- 0348
  X"c3",X"31",X"04",X"21",X"40",X"01",X"39",X"e5", -- 0350
  X"21",X"a6",X"04",X"e5",X"3e",X"02",X"cd",X"54", -- 0358
  X"17",X"c1",X"c1",X"7c",X"b5",X"c2",X"a9",X"03", -- 0360
  X"21",X"50",X"00",X"39",X"e5",X"3e",X"01",X"cd", -- 0368
  X"07",X"16",X"c1",X"7c",X"b5",X"ca",X"8d",X"03", -- 0370
  X"21",X"50",X"00",X"39",X"e5",X"3e",X"01",X"cd", -- 0378
  X"22",X"1b",X"c1",X"e5",X"3e",X"01",X"cd",X"33", -- 0380
  X"1f",X"c1",X"c3",X"a6",X"03",X"21",X"ab",X"04", -- 0388
  X"e5",X"3e",X"01",X"cd",X"ef",X"1d",X"c1",X"21", -- 0390
  X"50",X"00",X"39",X"e5",X"3e",X"01",X"cd",X"ef", -- 0398
  X"1d",X"c1",X"af",X"cd",X"5c",X"1c",X"c3",X"31", -- 03a0
  X"04",X"21",X"40",X"01",X"39",X"e5",X"21",X"b2", -- 03a8
  X"04",X"e5",X"3e",X"02",X"cd",X"54",X"17",X"c1", -- 03b0
  X"c1",X"7c",X"b5",X"c2",X"de",X"03",X"21",X"e2", -- 03b8
  X"01",X"39",X"e5",X"21",X"e4",X"01",X"39",X"cd", -- 03c0
  X"d5",X"27",X"e5",X"21",X"a4",X"00",X"39",X"e5", -- 03c8
  X"3e",X"02",X"cd",X"f4",X"08",X"c1",X"c1",X"d1", -- 03d0
  X"cd",X"15",X"28",X"c3",X"31",X"04",X"21",X"40", -- 03d8
  X"01",X"39",X"e5",X"3e",X"01",X"cd",X"07",X"16", -- 03e0
  X"c1",X"7c",X"b5",X"ca",X"05",X"04",X"21",X"e2", -- 03e8
  X"01",X"39",X"e5",X"21",X"42",X"01",X"39",X"e5", -- 03f0
  X"3e",X"01",X"cd",X"22",X"1b",X"c1",X"d1",X"cd", -- 03f8
  X"15",X"28",X"c3",X"31",X"04",X"21",X"e2",X"01", -- 0400
  X"39",X"e5",X"21",X"e4",X"01",X"39",X"cd",X"d5", -- 0408
  X"27",X"e5",X"21",X"44",X"01",X"39",X"e5",X"21", -- 0410
  X"56",X"00",X"39",X"e5",X"21",X"08",X"00",X"39", -- 0418
  X"e5",X"3e",X"04",X"cd",X"55",X"0e",X"eb",X"21", -- 0420
  X"08",X"00",X"39",X"f9",X"eb",X"d1",X"cd",X"15", -- 0428
  X"28",X"c3",X"73",X"01",X"21",X"e4",X"01",X"39", -- 0430
  X"f9",X"c9",X"4d",X"4f",X"4e",X"38",X"30",X"20", -- 0438
  X"56",X"65",X"72",X"73",X"69",X"6f",X"6e",X"20", -- 0440
  X"32",X"2e",X"32",X"20",X"53",X"42",X"43",X"38", -- 0448
  X"30",X"38",X"30",X"20",X"45",X"64",X"69",X"74", -- 0450
  X"69",X"6f",X"6e",X"00",X"49",X"6e",X"74",X"65", -- 0458
  X"6c",X"38",X"30",X"38",X"30",X"20",X"4d",X"6f", -- 0460
  X"6e",X"69",X"74",X"6f",X"72",X"20",X"50",X"72", -- 0468
  X"6f",X"67",X"72",X"61",X"6d",X"00",X"28",X"43", -- 0470
  X"29",X"31",X"39",X"39",X"36",X"2d",X"32",X"30", -- 0478
  X"31",X"38",X"20",X"4f",X"66",X"66",X"69",X"63", -- 0480
  X"65",X"20",X"54",X"45",X"54",X"53",X"55",X"00", -- 0488
  X"4c",X"49",X"53",X"54",X"00",X"44",X"55",X"4d", -- 0490
  X"50",X"00",X"53",X"59",X"53",X"54",X"45",X"4d", -- 0498
  X"00",X"48",X"45",X"4c",X"50",X"00",X"45",X"58", -- 04a0
  X"45",X"43",X"00",X"45",X"52",X"52",X"4f",X"52", -- 04a8
  X"2d",X"00",X"44",X"45",X"46",X"49",X"4e",X"45", -- 04b0
  X"00",X"21",X"04",X"00",X"39",X"e5",X"21",X"06", -- 04b8
  X"00",X"39",X"cd",X"d5",X"27",X"e5",X"3e",X"01", -- 04c0
  X"cd",X"ef",X"04",X"c1",X"d1",X"cd",X"15",X"28", -- 04c8
  X"21",X"04",X"00",X"39",X"cd",X"d5",X"27",X"eb", -- 04d0
  X"c1",X"e1",X"e5",X"c5",X"cd",X"7a",X"28",X"7c", -- 04d8
  X"b5",X"ca",X"e7",X"04",X"c3",X"b9",X"04",X"21", -- 04e0
  X"04",X"00",X"39",X"cd",X"d5",X"27",X"c9",X"3b", -- 04e8
  X"c5",X"21",X"20",X"00",X"e5",X"3e",X"01",X"cd", -- 04f0
  X"3e",X"1f",X"c1",X"21",X"05",X"00",X"39",X"cd", -- 04f8
  X"d5",X"27",X"e5",X"3e",X"01",X"cd",X"6a",X"1c", -- 0500
  X"c1",X"21",X"20",X"00",X"e5",X"3e",X"01",X"cd", -- 0508
  X"3e",X"1f",X"c1",X"21",X"02",X"00",X"39",X"e5", -- 0510
  X"21",X"07",X"00",X"39",X"54",X"5d",X"cd",X"d5", -- 0518
  X"27",X"23",X"cd",X"15",X"28",X"2b",X"cd",X"c8", -- 0520
  X"27",X"d1",X"7d",X"12",X"21",X"02",X"00",X"39", -- 0528
  X"cd",X"c8",X"27",X"e5",X"3e",X"01",X"cd",X"e0", -- 0530
  X"26",X"c1",X"e5",X"3e",X"01",X"cd",X"ef",X"1d", -- 0538
  X"c1",X"21",X"00",X"00",X"39",X"eb",X"21",X"05", -- 0540
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"15",X"28", -- 0548
  X"21",X"02",X"00",X"39",X"cd",X"c8",X"27",X"e5", -- 0550
  X"3e",X"01",X"cd",X"f1",X"26",X"c1",X"cd",X"d5", -- 0558
  X"27",X"eb",X"21",X"01",X"00",X"cd",X"30",X"28", -- 0560
  X"7c",X"b5",X"ca",X"9b",X"05",X"21",X"09",X"00", -- 0568
  X"e5",X"3e",X"01",X"cd",X"3e",X"1f",X"c1",X"21", -- 0570
  X"05",X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8", -- 0578
  X"27",X"e5",X"3e",X"01",X"cd",X"2f",X"1d",X"c1", -- 0580
  X"21",X"05",X"00",X"39",X"e5",X"cd",X"d5",X"27", -- 0588
  X"11",X"01",X"00",X"19",X"d1",X"cd",X"15",X"28", -- 0590
  X"c3",X"27",X"06",X"21",X"02",X"00",X"39",X"cd", -- 0598
  X"c8",X"27",X"e5",X"3e",X"01",X"cd",X"f1",X"26", -- 05a0
  X"c1",X"cd",X"d5",X"27",X"eb",X"21",X"02",X"00", -- 05a8
  X"cd",X"30",X"28",X"7c",X"b5",X"ca",X"e1",X"05", -- 05b0
  X"21",X"09",X"00",X"e5",X"3e",X"01",X"cd",X"3e", -- 05b8
  X"1f",X"c1",X"e1",X"e5",X"cd",X"d5",X"27",X"e5", -- 05c0
  X"3e",X"01",X"cd",X"6a",X"1c",X"c1",X"21",X"05", -- 05c8
  X"00",X"39",X"e5",X"cd",X"d5",X"27",X"11",X"02", -- 05d0
  X"00",X"19",X"d1",X"cd",X"15",X"28",X"c3",X"27", -- 05d8
  X"06",X"21",X"02",X"00",X"39",X"cd",X"c8",X"27", -- 05e0
  X"e5",X"3e",X"01",X"cd",X"f1",X"26",X"c1",X"cd", -- 05e8
  X"d5",X"27",X"7c",X"b5",X"ca",X"19",X"06",X"21", -- 05f0
  X"09",X"00",X"e5",X"3e",X"01",X"cd",X"3e",X"1f", -- 05f8
  X"c1",X"21",X"02",X"00",X"39",X"cd",X"c8",X"27", -- 0600
  X"e5",X"3e",X"01",X"cd",X"f1",X"26",X"c1",X"e5", -- 0608
  X"3e",X"01",X"cd",X"ef",X"1d",X"c1",X"c3",X"27", -- 0610
  X"06",X"af",X"cd",X"5c",X"1c",X"21",X"05",X"00", -- 0618
  X"39",X"cd",X"d5",X"27",X"33",X"c1",X"c9",X"21", -- 0620
  X"00",X"00",X"39",X"eb",X"21",X"05",X"00",X"39", -- 0628
  X"cd",X"d5",X"27",X"cd",X"15",X"28",X"21",X"02", -- 0630
  X"00",X"39",X"cd",X"c8",X"27",X"e5",X"3e",X"01", -- 0638
  X"cd",X"02",X"27",X"c1",X"cd",X"d5",X"27",X"eb", -- 0640
  X"21",X"01",X"00",X"cd",X"30",X"28",X"7c",X"b5", -- 0648
  X"ca",X"81",X"06",X"21",X"2c",X"00",X"e5",X"3e", -- 0650
  X"01",X"cd",X"3e",X"1f",X"c1",X"21",X"05",X"00", -- 0658
  X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"e5", -- 0660
  X"3e",X"01",X"cd",X"2f",X"1d",X"c1",X"21",X"05", -- 0668
  X"00",X"39",X"e5",X"cd",X"d5",X"27",X"11",X"01", -- 0670
  X"00",X"19",X"d1",X"cd",X"15",X"28",X"c3",X"fc", -- 0678
  X"06",X"21",X"02",X"00",X"39",X"cd",X"c8",X"27", -- 0680
  X"e5",X"3e",X"01",X"cd",X"02",X"27",X"c1",X"cd", -- 0688
  X"d5",X"27",X"eb",X"21",X"02",X"00",X"cd",X"30", -- 0690
  X"28",X"7c",X"b5",X"ca",X"c7",X"06",X"21",X"2c", -- 0698
  X"00",X"e5",X"3e",X"01",X"cd",X"3e",X"1f",X"c1", -- 06a0
  X"e1",X"e5",X"cd",X"d5",X"27",X"e5",X"3e",X"01", -- 06a8
  X"cd",X"6a",X"1c",X"c1",X"21",X"05",X"00",X"39", -- 06b0
  X"e5",X"cd",X"d5",X"27",X"11",X"02",X"00",X"19", -- 06b8
  X"d1",X"cd",X"15",X"28",X"c3",X"fc",X"06",X"21", -- 06c0
  X"02",X"00",X"39",X"cd",X"c8",X"27",X"e5",X"3e", -- 06c8
  X"01",X"cd",X"02",X"27",X"c1",X"cd",X"d5",X"27", -- 06d0
  X"7c",X"b5",X"ca",X"fc",X"06",X"21",X"2c",X"00", -- 06d8
  X"e5",X"3e",X"01",X"cd",X"3e",X"1f",X"c1",X"21", -- 06e0
  X"02",X"00",X"39",X"cd",X"c8",X"27",X"e5",X"3e", -- 06e8
  X"01",X"cd",X"02",X"27",X"c1",X"e5",X"3e",X"01", -- 06f0
  X"cd",X"ef",X"1d",X"c1",X"af",X"cd",X"5c",X"1c", -- 06f8
  X"21",X"05",X"00",X"39",X"cd",X"d5",X"27",X"33", -- 0700
  X"c1",X"c9",X"21",X"80",X"07",X"e5",X"3e",X"01", -- 0708
  X"cd",X"ef",X"1d",X"c1",X"21",X"87",X"07",X"e5", -- 0710
  X"3e",X"01",X"cd",X"ef",X"1d",X"c1",X"21",X"b8", -- 0718
  X"07",X"e5",X"3e",X"01",X"cd",X"ef",X"1d",X"c1", -- 0720
  X"af",X"cd",X"5c",X"1c",X"21",X"04",X"00",X"39", -- 0728
  X"e5",X"21",X"06",X"00",X"39",X"cd",X"d5",X"27", -- 0730
  X"eb",X"21",X"f0",X"ff",X"cd",X"29",X"28",X"d1", -- 0738
  X"cd",X"15",X"28",X"21",X"04",X"00",X"39",X"e5", -- 0740
  X"21",X"06",X"00",X"39",X"cd",X"d5",X"27",X"e5", -- 0748
  X"3e",X"01",X"cd",X"be",X"07",X"c1",X"d1",X"cd", -- 0750
  X"15",X"28",X"21",X"04",X"00",X"39",X"cd",X"d5", -- 0758
  X"27",X"eb",X"21",X"01",X"00",X"cd",X"8c",X"28", -- 0760
  X"eb",X"c1",X"e1",X"e5",X"c5",X"cd",X"6d",X"28", -- 0768
  X"7c",X"b5",X"ca",X"78",X"07",X"c3",X"43",X"07", -- 0770
  X"21",X"04",X"00",X"39",X"cd",X"d5",X"27",X"c9", -- 0778
  X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"2b", -- 0780
  X"30",X"20",X"2b",X"31",X"20",X"2b",X"32",X"20", -- 0788
  X"2b",X"33",X"20",X"2b",X"34",X"20",X"2b",X"35", -- 0790
  X"20",X"2b",X"36",X"20",X"2b",X"37",X"20",X"2b", -- 0798
  X"38",X"20",X"2b",X"39",X"20",X"2b",X"41",X"20", -- 07a0
  X"2b",X"42",X"20",X"2b",X"43",X"20",X"2b",X"44", -- 07a8
  X"20",X"2b",X"45",X"20",X"2b",X"46",X"20",X"00", -- 07b0
  X"41",X"53",X"43",X"49",X"49",X"00",X"21",X"ee", -- 07b8
  X"ff",X"39",X"f9",X"21",X"20",X"00",X"e5",X"3e", -- 07c0
  X"01",X"cd",X"3e",X"1f",X"c1",X"21",X"14",X"00", -- 07c8
  X"39",X"cd",X"d5",X"27",X"e5",X"3e",X"01",X"cd", -- 07d0
  X"6a",X"1c",X"c1",X"21",X"20",X"00",X"e5",X"3e", -- 07d8
  X"01",X"cd",X"3e",X"1f",X"c1",X"21",X"00",X"00", -- 07e0
  X"39",X"eb",X"21",X"00",X"00",X"cd",X"15",X"28", -- 07e8
  X"d1",X"d5",X"21",X"10",X"00",X"cd",X"50",X"28", -- 07f0
  X"7c",X"b5",X"ca",X"31",X"08",X"c3",X"11",X"08", -- 07f8
  X"21",X"00",X"00",X"39",X"54",X"5d",X"cd",X"d5", -- 0800
  X"27",X"23",X"cd",X"15",X"28",X"2b",X"c3",X"f0", -- 0808
  X"07",X"21",X"02",X"00",X"39",X"eb",X"e1",X"e5", -- 0810
  X"19",X"e5",X"21",X"16",X"00",X"39",X"54",X"5d", -- 0818
  X"cd",X"d5",X"27",X"23",X"cd",X"15",X"28",X"2b", -- 0820
  X"cd",X"c8",X"27",X"d1",X"7d",X"12",X"c3",X"00", -- 0828
  X"08",X"21",X"00",X"00",X"39",X"eb",X"21",X"00", -- 0830
  X"00",X"cd",X"15",X"28",X"d1",X"d5",X"21",X"10", -- 0838
  X"00",X"cd",X"50",X"28",X"7c",X"b5",X"ca",X"7c", -- 0840
  X"08",X"c3",X"5d",X"08",X"21",X"00",X"00",X"39", -- 0848
  X"54",X"5d",X"cd",X"d5",X"27",X"23",X"cd",X"15", -- 0850
  X"28",X"2b",X"c3",X"3c",X"08",X"21",X"02",X"00", -- 0858
  X"39",X"eb",X"e1",X"e5",X"19",X"cd",X"c8",X"27", -- 0860
  X"e5",X"3e",X"01",X"cd",X"2f",X"1d",X"c1",X"21", -- 0868
  X"20",X"00",X"e5",X"3e",X"01",X"cd",X"3e",X"1f", -- 0870
  X"c1",X"c3",X"4c",X"08",X"21",X"00",X"00",X"39", -- 0878
  X"eb",X"21",X"00",X"00",X"cd",X"15",X"28",X"d1", -- 0880
  X"d5",X"21",X"10",X"00",X"cd",X"50",X"28",X"7c", -- 0888
  X"b5",X"ca",X"e1",X"08",X"c3",X"a8",X"08",X"21", -- 0890
  X"00",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 0898
  X"23",X"cd",X"15",X"28",X"2b",X"c3",X"87",X"08", -- 08a0
  X"21",X"02",X"00",X"39",X"eb",X"e1",X"e5",X"19", -- 08a8
  X"cd",X"c8",X"27",X"e5",X"3e",X"01",X"cd",X"bf", -- 08b0
  X"14",X"c1",X"7c",X"b5",X"ca",X"d4",X"08",X"21", -- 08b8
  X"02",X"00",X"39",X"eb",X"e1",X"e5",X"19",X"cd", -- 08c0
  X"c8",X"27",X"e5",X"3e",X"01",X"cd",X"3e",X"1f", -- 08c8
  X"c1",X"c3",X"de",X"08",X"21",X"2e",X"00",X"e5", -- 08d0
  X"3e",X"01",X"cd",X"3e",X"1f",X"c1",X"c3",X"97", -- 08d8
  X"08",X"af",X"cd",X"5c",X"1c",X"21",X"14",X"00", -- 08e0
  X"39",X"cd",X"d5",X"27",X"eb",X"21",X"12",X"00", -- 08e8
  X"39",X"f9",X"eb",X"c9",X"21",X"ae",X"ff",X"39", -- 08f0
  X"f9",X"21",X"54",X"00",X"39",X"cd",X"d5",X"27", -- 08f8
  X"cd",X"c8",X"27",X"7c",X"b5",X"ca",X"ef",X"09", -- 0900
  X"21",X"54",X"00",X"39",X"cd",X"d5",X"27",X"e5", -- 0908
  X"21",X"04",X"00",X"39",X"e5",X"21",X"58",X"00", -- 0910
  X"39",X"cd",X"d5",X"27",X"e5",X"3e",X"03",X"cd", -- 0918
  X"35",X"13",X"c1",X"c1",X"c1",X"21",X"00",X"00", -- 0920
  X"39",X"eb",X"21",X"02",X"00",X"39",X"cd",X"15", -- 0928
  X"28",X"e1",X"e5",X"e5",X"3e",X"01",X"cd",X"07", -- 0930
  X"16",X"c1",X"7c",X"b5",X"ca",X"5f",X"09",X"21", -- 0938
  X"56",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 0940
  X"23",X"cd",X"15",X"28",X"2b",X"e5",X"c1",X"e1", -- 0948
  X"e5",X"c5",X"e5",X"3e",X"01",X"cd",X"e9",X"19", -- 0950
  X"c1",X"d1",X"7d",X"12",X"c3",X"ec",X"09",X"e1", -- 0958
  X"e5",X"cd",X"c8",X"27",X"eb",X"21",X"27",X"00", -- 0960
  X"cd",X"30",X"28",X"7c",X"b5",X"ca",X"d0",X"09", -- 0968
  X"21",X"00",X"00",X"39",X"54",X"5d",X"cd",X"d5", -- 0970
  X"27",X"23",X"cd",X"15",X"28",X"2b",X"e1",X"e5", -- 0978
  X"cd",X"c8",X"27",X"7c",X"b5",X"ca",X"9f",X"09", -- 0980
  X"e1",X"e5",X"cd",X"c8",X"27",X"eb",X"21",X"27", -- 0988
  X"00",X"cd",X"36",X"28",X"7c",X"b5",X"ca",X"9f", -- 0990
  X"09",X"21",X"01",X"00",X"c3",X"a2",X"09",X"21", -- 0998
  X"00",X"00",X"7c",X"b5",X"ca",X"cd",X"09",X"21", -- 09a0
  X"56",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 09a8
  X"23",X"cd",X"15",X"28",X"2b",X"e5",X"21",X"02", -- 09b0
  X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27",X"23", -- 09b8
  X"cd",X"15",X"28",X"2b",X"cd",X"c8",X"27",X"d1", -- 09c0
  X"7d",X"12",X"c3",X"7e",X"09",X"c3",X"ec",X"09", -- 09c8
  X"21",X"fe",X"09",X"e5",X"3e",X"01",X"cd",X"ef", -- 09d0
  X"1d",X"c1",X"21",X"02",X"00",X"39",X"e5",X"3e", -- 09d8
  X"01",X"cd",X"ef",X"1d",X"c1",X"af",X"cd",X"5c", -- 09e0
  X"1c",X"c3",X"ef",X"09",X"c3",X"f9",X"08",X"21", -- 09e8
  X"56",X"00",X"39",X"cd",X"d5",X"27",X"eb",X"21", -- 09f0
  X"52",X"00",X"39",X"f9",X"eb",X"c9",X"45",X"72", -- 09f8
  X"72",X"6f",X"72",X"2d",X"00",X"c5",X"c5",X"c5", -- 0a00
  X"21",X"08",X"00",X"39",X"cd",X"d5",X"27",X"cd", -- 0a08
  X"c8",X"27",X"7c",X"b5",X"c2",X"8a",X"0a",X"21", -- 0a10
  X"4c",X"0d",X"e5",X"3e",X"01",X"cd",X"ef",X"1d", -- 0a18
  X"c1",X"af",X"cd",X"5c",X"1c",X"21",X"72",X"0d", -- 0a20
  X"e5",X"3e",X"01",X"cd",X"ef",X"1d",X"c1",X"af", -- 0a28
  X"cd",X"5c",X"1c",X"21",X"8a",X"0d",X"e5",X"3e", -- 0a30
  X"01",X"cd",X"ef",X"1d",X"c1",X"af",X"cd",X"5c", -- 0a38
  X"1c",X"21",X"a5",X"0d",X"e5",X"3e",X"01",X"cd", -- 0a40
  X"ef",X"1d",X"c1",X"af",X"cd",X"5c",X"1c",X"21", -- 0a48
  X"c0",X"0d",X"e5",X"3e",X"01",X"cd",X"ef",X"1d", -- 0a50
  X"c1",X"af",X"cd",X"5c",X"1c",X"21",X"dc",X"0d", -- 0a58
  X"e5",X"3e",X"01",X"cd",X"ef",X"1d",X"c1",X"af", -- 0a60
  X"cd",X"5c",X"1c",X"21",X"fb",X"0d",X"e5",X"3e", -- 0a68
  X"01",X"cd",X"ef",X"1d",X"c1",X"af",X"cd",X"5c", -- 0a70
  X"1c",X"21",X"17",X"0e",X"e5",X"3e",X"01",X"cd", -- 0a78
  X"ef",X"1d",X"c1",X"af",X"cd",X"5c",X"1c",X"c3", -- 0a80
  X"48",X"0d",X"21",X"08",X"00",X"39",X"cd",X"d5", -- 0a88
  X"27",X"cd",X"c8",X"27",X"eb",X"21",X"00",X"00", -- 0a90
  X"cd",X"36",X"28",X"7c",X"b5",X"ca",X"e0",X"0a", -- 0a98
  X"21",X"08",X"00",X"39",X"cd",X"d5",X"27",X"cd", -- 0aa0
  X"c8",X"27",X"e5",X"3e",X"01",X"cd",X"ef",X"14", -- 0aa8
  X"c1",X"7c",X"b5",X"c2",X"d2",X"0a",X"21",X"08", -- 0ab0
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27", -- 0ab8
  X"eb",X"21",X"2c",X"00",X"cd",X"30",X"28",X"7c", -- 0ac0
  X"b5",X"c2",X"d2",X"0a",X"21",X"00",X"00",X"c3", -- 0ac8
  X"d5",X"0a",X"21",X"01",X"00",X"7c",X"b5",X"ca", -- 0ad0
  X"e0",X"0a",X"21",X"01",X"00",X"c3",X"e3",X"0a", -- 0ad8
  X"21",X"00",X"00",X"7c",X"b5",X"ca",X"f9",X"0a", -- 0ae0
  X"21",X"08",X"00",X"39",X"54",X"5d",X"cd",X"d5", -- 0ae8
  X"27",X"23",X"cd",X"15",X"28",X"2b",X"c3",X"8a", -- 0af0
  X"0a",X"21",X"04",X"00",X"39",X"eb",X"21",X"08", -- 0af8
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"15",X"28", -- 0b00
  X"21",X"04",X"00",X"39",X"cd",X"d5",X"27",X"cd", -- 0b08
  X"c8",X"27",X"eb",X"21",X"00",X"00",X"cd",X"36", -- 0b10
  X"28",X"7c",X"b5",X"ca",X"53",X"0b",X"21",X"04", -- 0b18
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27", -- 0b20
  X"e5",X"3e",X"01",X"cd",X"ef",X"14",X"c1",X"cd", -- 0b28
  X"9f",X"28",X"7c",X"b5",X"ca",X"53",X"0b",X"21", -- 0b30
  X"04",X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8", -- 0b38
  X"27",X"eb",X"21",X"2c",X"00",X"cd",X"36",X"28", -- 0b40
  X"7c",X"b5",X"ca",X"53",X"0b",X"21",X"01",X"00", -- 0b48
  X"c3",X"56",X"0b",X"21",X"00",X"00",X"7c",X"b5", -- 0b50
  X"ca",X"6c",X"0b",X"21",X"04",X"00",X"39",X"54", -- 0b58
  X"5d",X"cd",X"d5",X"27",X"23",X"cd",X"15",X"28", -- 0b60
  X"2b",X"c3",X"08",X"0b",X"21",X"04",X"00",X"39", -- 0b68
  X"cd",X"d5",X"27",X"eb",X"21",X"00",X"00",X"7d", -- 0b70
  X"12",X"21",X"00",X"00",X"39",X"eb",X"21",X"00", -- 0b78
  X"00",X"cd",X"15",X"28",X"21",X"02",X"00",X"39", -- 0b80
  X"eb",X"21",X"00",X"00",X"cd",X"15",X"28",X"c1", -- 0b88
  X"d1",X"d5",X"c5",X"21",X"ff",X"00",X"cd",X"43", -- 0b90
  X"28",X"7c",X"b5",X"ca",X"25",X"0d",X"c3",X"b2", -- 0b98
  X"0b",X"21",X"02",X"00",X"39",X"54",X"5d",X"cd", -- 0ba0
  X"d5",X"27",X"23",X"cd",X"15",X"28",X"2b",X"c3", -- 0ba8
  X"8f",X"0b",X"21",X"08",X"00",X"39",X"cd",X"d5", -- 0bb0
  X"27",X"e5",X"21",X"04",X"00",X"39",X"cd",X"d5", -- 0bb8
  X"27",X"e5",X"3e",X"01",X"cd",X"e0",X"26",X"c1", -- 0bc0
  X"e5",X"3e",X"02",X"cd",X"54",X"17",X"c1",X"c1", -- 0bc8
  X"7c",X"b5",X"c2",X"22",X"0d",X"21",X"37",X"0e", -- 0bd0
  X"e5",X"3e",X"01",X"cd",X"ef",X"1d",X"c1",X"c1", -- 0bd8
  X"e1",X"e5",X"c5",X"e5",X"3e",X"01",X"cd",X"e0", -- 0be0
  X"26",X"c1",X"e5",X"3e",X"01",X"cd",X"ef",X"1d", -- 0be8
  X"c1",X"c1",X"e1",X"e5",X"c5",X"e5",X"3e",X"01", -- 0bf0
  X"cd",X"f1",X"26",X"c1",X"cd",X"d5",X"27",X"eb", -- 0bf8
  X"21",X"01",X"00",X"cd",X"30",X"28",X"7c",X"b5", -- 0c00
  X"ca",X"22",X"0c",X"21",X"09",X"00",X"e5",X"3e", -- 0c08
  X"01",X"cd",X"3e",X"1f",X"c1",X"21",X"3e",X"0e", -- 0c10
  X"e5",X"3e",X"01",X"cd",X"ef",X"1d",X"c1",X"c3", -- 0c18
  X"82",X"0c",X"c1",X"e1",X"e5",X"c5",X"e5",X"3e", -- 0c20
  X"01",X"cd",X"f1",X"26",X"c1",X"cd",X"d5",X"27", -- 0c28
  X"eb",X"21",X"02",X"00",X"cd",X"30",X"28",X"7c", -- 0c30
  X"b5",X"ca",X"53",X"0c",X"21",X"09",X"00",X"e5", -- 0c38
  X"3e",X"01",X"cd",X"3e",X"1f",X"c1",X"21",X"41", -- 0c40
  X"0e",X"e5",X"3e",X"01",X"cd",X"ef",X"1d",X"c1", -- 0c48
  X"c3",X"82",X"0c",X"c1",X"e1",X"e5",X"c5",X"e5", -- 0c50
  X"3e",X"01",X"cd",X"f1",X"26",X"c1",X"cd",X"d5", -- 0c58
  X"27",X"7c",X"b5",X"ca",X"82",X"0c",X"21",X"09", -- 0c60
  X"00",X"e5",X"3e",X"01",X"cd",X"3e",X"1f",X"c1", -- 0c68
  X"c1",X"e1",X"e5",X"c5",X"e5",X"3e",X"01",X"cd", -- 0c70
  X"f1",X"26",X"c1",X"e5",X"3e",X"01",X"cd",X"ef", -- 0c78
  X"1d",X"c1",X"c1",X"e1",X"e5",X"c5",X"e5",X"3e", -- 0c80
  X"01",X"cd",X"02",X"27",X"c1",X"cd",X"d5",X"27", -- 0c88
  X"eb",X"21",X"01",X"00",X"cd",X"30",X"28",X"7c", -- 0c90
  X"b5",X"ca",X"b3",X"0c",X"21",X"2c",X"00",X"e5", -- 0c98
  X"3e",X"01",X"cd",X"3e",X"1f",X"c1",X"21",X"46", -- 0ca0
  X"0e",X"e5",X"3e",X"01",X"cd",X"ef",X"1d",X"c1", -- 0ca8
  X"c3",X"13",X"0d",X"c1",X"e1",X"e5",X"c5",X"e5", -- 0cb0
  X"3e",X"01",X"cd",X"02",X"27",X"c1",X"cd",X"d5", -- 0cb8
  X"27",X"eb",X"21",X"02",X"00",X"cd",X"30",X"28", -- 0cc0
  X"7c",X"b5",X"ca",X"e4",X"0c",X"21",X"2c",X"00", -- 0cc8
  X"e5",X"3e",X"01",X"cd",X"3e",X"1f",X"c1",X"21", -- 0cd0
  X"49",X"0e",X"e5",X"3e",X"01",X"cd",X"ef",X"1d", -- 0cd8
  X"c1",X"c3",X"13",X"0d",X"c1",X"e1",X"e5",X"c5", -- 0ce0
  X"e5",X"3e",X"01",X"cd",X"02",X"27",X"c1",X"cd", -- 0ce8
  X"d5",X"27",X"7c",X"b5",X"ca",X"13",X"0d",X"21", -- 0cf0
  X"2c",X"00",X"e5",X"3e",X"01",X"cd",X"3e",X"1f", -- 0cf8
  X"c1",X"c1",X"e1",X"e5",X"c5",X"e5",X"3e",X"01", -- 0d00
  X"cd",X"02",X"27",X"c1",X"e5",X"3e",X"01",X"cd", -- 0d08
  X"ef",X"1d",X"c1",X"af",X"cd",X"5c",X"1c",X"21", -- 0d10
  X"00",X"00",X"39",X"eb",X"21",X"01",X"00",X"cd", -- 0d18
  X"15",X"28",X"c3",X"a1",X"0b",X"e1",X"e5",X"7c", -- 0d20
  X"b5",X"c2",X"48",X"0d",X"21",X"4e",X"0e",X"e5", -- 0d28
  X"3e",X"01",X"cd",X"ef",X"1d",X"c1",X"21",X"08", -- 0d30
  X"00",X"39",X"cd",X"d5",X"27",X"e5",X"3e",X"01", -- 0d38
  X"cd",X"ef",X"1d",X"c1",X"af",X"cd",X"5c",X"1c", -- 0d40
  X"c1",X"c1",X"c1",X"c9",X"20",X"20",X"20",X"20", -- 0d48
  X"20",X"20",X"78",X"78",X"78",X"78",X"20",X"20", -- 0d50
  X"20",X"20",X"20",X"43",X"68",X"61",X"6e",X"67", -- 0d58
  X"65",X"20",X"63",X"75",X"72",X"72",X"65",X"6e", -- 0d60
  X"74",X"20",X"61",X"64",X"64",X"72",X"65",X"73", -- 0d68
  X"73",X"00",X"20",X"20",X"20",X"20",X"20",X"20", -- 0d70
  X"6d",X"6e",X"65",X"6d",X"6f",X"6e",X"69",X"63", -- 0d78
  X"20",X"41",X"73",X"73",X"65",X"6d",X"62",X"6c", -- 0d80
  X"65",X"00",X"20",X"20",X"20",X"20",X"20",X"20", -- 0d88
  X"4c",X"49",X"53",X"54",X"20",X"20",X"20",X"20", -- 0d90
  X"20",X"44",X"69",X"73",X"61",X"73",X"73",X"65", -- 0d98
  X"6d",X"62",X"6c",X"65",X"00",X"20",X"20",X"20", -- 0da0
  X"20",X"20",X"20",X"44",X"45",X"46",X"49",X"4e", -- 0da8
  X"45",X"20",X"20",X"20",X"44",X"65",X"66",X"69", -- 0db0
  X"6e",X"65",X"20",X"64",X"61",X"74",X"61",X"00", -- 0db8
  X"20",X"20",X"20",X"20",X"20",X"20",X"44",X"55", -- 0dc0
  X"4d",X"50",X"20",X"20",X"20",X"20",X"20",X"44", -- 0dc8
  X"69",X"73",X"70",X"6c",X"61",X"79",X"20",X"64", -- 0dd0
  X"61",X"74",X"61",X"00",X"20",X"20",X"20",X"20", -- 0dd8
  X"20",X"20",X"45",X"58",X"45",X"43",X"20",X"20", -- 0de0
  X"20",X"20",X"20",X"45",X"78",X"65",X"63",X"75", -- 0de8
  X"74",X"65",X"20",X"70",X"72",X"6f",X"67",X"72", -- 0df0
  X"61",X"6d",X"00",X"20",X"20",X"20",X"20",X"20", -- 0df8
  X"20",X"48",X"45",X"4c",X"50",X"20",X"20",X"20", -- 0e00
  X"20",X"20",X"44",X"69",X"73",X"70",X"6c",X"61", -- 0e08
  X"79",X"20",X"68",X"65",X"6c",X"70",X"00",X"20", -- 0e10
  X"20",X"20",X"20",X"20",X"20",X"53",X"59",X"53", -- 0e18
  X"54",X"45",X"4d",X"20",X"20",X"20",X"52",X"65", -- 0e20
  X"74",X"75",X"72",X"6e",X"20",X"74",X"6f",X"20", -- 0e28
  X"73",X"79",X"73",X"74",X"65",X"6d",X"00",X"20", -- 0e30
  X"20",X"20",X"20",X"20",X"20",X"00",X"78",X"78", -- 0e38
  X"00",X"78",X"78",X"78",X"78",X"00",X"78",X"78", -- 0e40
  X"00",X"78",X"78",X"78",X"78",X"00",X"45",X"52", -- 0e48
  X"52",X"4f",X"52",X"2d",X"00",X"3b",X"c5",X"c5", -- 0e50
  X"21",X"04",X"00",X"39",X"eb",X"21",X"ff",X"00", -- 0e58
  X"7d",X"12",X"21",X"00",X"00",X"39",X"eb",X"21", -- 0e60
  X"00",X"00",X"cd",X"15",X"28",X"21",X"04",X"00", -- 0e68
  X"39",X"54",X"5d",X"cd",X"c8",X"27",X"2b",X"7d", -- 0e70
  X"12",X"23",X"7c",X"b5",X"ca",X"92",X"0e",X"d1", -- 0e78
  X"d5",X"21",X"00",X"00",X"cd",X"30",X"28",X"7c", -- 0e80
  X"b5",X"ca",X"92",X"0e",X"21",X"01",X"00",X"c3", -- 0e88
  X"95",X"0e",X"21",X"00",X"00",X"7c",X"b5",X"ca", -- 0e90
  X"b7",X"0f",X"21",X"0b",X"00",X"39",X"cd",X"d5", -- 0e98
  X"27",X"e5",X"21",X"06",X"00",X"39",X"cd",X"c8", -- 0ea0
  X"27",X"e5",X"3e",X"01",X"cd",X"e0",X"26",X"c1", -- 0ea8
  X"e5",X"3e",X"02",X"cd",X"54",X"17",X"c1",X"c1", -- 0eb0
  X"7c",X"b5",X"c2",X"b4",X"0f",X"21",X"09",X"00", -- 0eb8
  X"39",X"cd",X"d5",X"27",X"e5",X"21",X"06",X"00", -- 0ec0
  X"39",X"cd",X"c8",X"27",X"e5",X"3e",X"01",X"cd", -- 0ec8
  X"f1",X"26",X"c1",X"e5",X"3e",X"02",X"cd",X"54", -- 0ed0
  X"17",X"c1",X"c1",X"eb",X"21",X"00",X"00",X"cd", -- 0ed8
  X"30",X"28",X"7c",X"b5",X"c2",X"2b",X"0f",X"21", -- 0ee0
  X"09",X"00",X"39",X"cd",X"d5",X"27",X"e5",X"3e", -- 0ee8
  X"01",X"cd",X"07",X"16",X"c1",X"7c",X"b5",X"ca", -- 0ef0
  X"1d",X"0f",X"21",X"04",X"00",X"39",X"cd",X"c8", -- 0ef8
  X"27",X"e5",X"3e",X"01",X"cd",X"f1",X"26",X"c1", -- 0f00
  X"cd",X"d5",X"27",X"eb",X"21",X"02",X"00",X"cd", -- 0f08
  X"43",X"28",X"7c",X"b5",X"ca",X"1d",X"0f",X"21", -- 0f10
  X"01",X"00",X"c3",X"20",X"0f",X"21",X"00",X"00", -- 0f18
  X"7c",X"b5",X"c2",X"2b",X"0f",X"21",X"00",X"00", -- 0f20
  X"c3",X"2e",X"0f",X"21",X"01",X"00",X"7c",X"b5", -- 0f28
  X"ca",X"b4",X"0f",X"21",X"07",X"00",X"39",X"cd", -- 0f30
  X"d5",X"27",X"e5",X"21",X"06",X"00",X"39",X"cd", -- 0f38
  X"c8",X"27",X"e5",X"3e",X"01",X"cd",X"02",X"27", -- 0f40
  X"c1",X"e5",X"3e",X"02",X"cd",X"54",X"17",X"c1", -- 0f48
  X"c1",X"eb",X"21",X"00",X"00",X"cd",X"30",X"28", -- 0f50
  X"7c",X"b5",X"c2",X"a1",X"0f",X"21",X"07",X"00", -- 0f58
  X"39",X"cd",X"d5",X"27",X"e5",X"3e",X"01",X"cd", -- 0f60
  X"07",X"16",X"c1",X"7c",X"b5",X"ca",X"93",X"0f", -- 0f68
  X"21",X"04",X"00",X"39",X"cd",X"c8",X"27",X"e5", -- 0f70
  X"3e",X"01",X"cd",X"02",X"27",X"c1",X"cd",X"d5", -- 0f78
  X"27",X"eb",X"21",X"02",X"00",X"cd",X"43",X"28", -- 0f80
  X"7c",X"b5",X"ca",X"93",X"0f",X"21",X"01",X"00", -- 0f88
  X"c3",X"96",X"0f",X"21",X"00",X"00",X"7c",X"b5", -- 0f90
  X"c2",X"a1",X"0f",X"21",X"00",X"00",X"c3",X"a4", -- 0f98
  X"0f",X"21",X"01",X"00",X"7c",X"b5",X"ca",X"b4", -- 0fa0
  X"0f",X"21",X"00",X"00",X"39",X"eb",X"21",X"01", -- 0fa8
  X"00",X"cd",X"15",X"28",X"c3",X"6d",X"0e",X"e1", -- 0fb0
  X"e5",X"7c",X"b5",X"c2",X"33",X"10",X"21",X"8f", -- 0fb8
  X"11",X"e5",X"3e",X"01",X"cd",X"ef",X"1d",X"c1", -- 0fc0
  X"21",X"0b",X"00",X"39",X"cd",X"d5",X"27",X"e5", -- 0fc8
  X"3e",X"01",X"cd",X"ef",X"1d",X"c1",X"21",X"20", -- 0fd0
  X"00",X"e5",X"3e",X"01",X"cd",X"3e",X"1f",X"c1", -- 0fd8
  X"21",X"09",X"00",X"39",X"cd",X"d5",X"27",X"cd", -- 0fe0
  X"c8",X"27",X"7c",X"b5",X"ca",X"fd",X"0f",X"21", -- 0fe8
  X"09",X"00",X"39",X"cd",X"d5",X"27",X"e5",X"3e", -- 0ff0
  X"01",X"cd",X"ef",X"1d",X"c1",X"21",X"07",X"00", -- 0ff8
  X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"7c", -- 1000
  X"b5",X"ca",X"24",X"10",X"21",X"2c",X"00",X"e5", -- 1008
  X"3e",X"01",X"cd",X"3e",X"1f",X"c1",X"21",X"07", -- 1010
  X"00",X"39",X"cd",X"d5",X"27",X"e5",X"3e",X"01", -- 1018
  X"cd",X"ef",X"1d",X"c1",X"af",X"cd",X"5c",X"1c", -- 1020
  X"21",X"0d",X"00",X"39",X"cd",X"d5",X"27",X"33", -- 1028
  X"c1",X"c1",X"c9",X"21",X"04",X"00",X"39",X"54", -- 1030
  X"5d",X"cd",X"c8",X"27",X"23",X"7d",X"12",X"2b", -- 1038
  X"21",X"0d",X"00",X"39",X"54",X"5d",X"cd",X"d5", -- 1040
  X"27",X"23",X"cd",X"15",X"28",X"2b",X"eb",X"21", -- 1048
  X"04",X"00",X"39",X"cd",X"c8",X"27",X"7d",X"12", -- 1050
  X"21",X"02",X"00",X"39",X"eb",X"21",X"0d",X"00", -- 1058
  X"39",X"cd",X"d5",X"27",X"cd",X"15",X"28",X"21", -- 1060
  X"04",X"00",X"39",X"cd",X"c8",X"27",X"e5",X"3e", -- 1068
  X"01",X"cd",X"f1",X"26",X"c1",X"cd",X"d5",X"27", -- 1070
  X"eb",X"21",X"01",X"00",X"cd",X"30",X"28",X"7c", -- 1078
  X"b5",X"ca",X"b0",X"10",X"21",X"0d",X"00",X"39", -- 1080
  X"cd",X"d5",X"27",X"e5",X"21",X"0b",X"00",X"39", -- 1088
  X"cd",X"d5",X"27",X"e5",X"3e",X"01",X"cd",X"e9", -- 1090
  X"19",X"c1",X"d1",X"7d",X"12",X"21",X"0d",X"00", -- 1098
  X"39",X"e5",X"cd",X"d5",X"27",X"11",X"01",X"00", -- 10a0
  X"19",X"d1",X"cd",X"15",X"28",X"c3",X"84",X"11", -- 10a8
  X"21",X"04",X"00",X"39",X"cd",X"c8",X"27",X"e5", -- 10b0
  X"3e",X"01",X"cd",X"02",X"27",X"c1",X"cd",X"d5", -- 10b8
  X"27",X"eb",X"21",X"01",X"00",X"cd",X"30",X"28", -- 10c0
  X"7c",X"b5",X"ca",X"f9",X"10",X"21",X"0d",X"00", -- 10c8
  X"39",X"cd",X"d5",X"27",X"e5",X"21",X"09",X"00", -- 10d0
  X"39",X"cd",X"d5",X"27",X"e5",X"3e",X"01",X"cd", -- 10d8
  X"e9",X"19",X"c1",X"d1",X"7d",X"12",X"21",X"0d", -- 10e0
  X"00",X"39",X"e5",X"cd",X"d5",X"27",X"11",X"01", -- 10e8
  X"00",X"19",X"d1",X"cd",X"15",X"28",X"c3",X"84", -- 10f0
  X"11",X"21",X"04",X"00",X"39",X"cd",X"c8",X"27", -- 10f8
  X"e5",X"3e",X"01",X"cd",X"f1",X"26",X"c1",X"cd", -- 1100
  X"d5",X"27",X"eb",X"21",X"02",X"00",X"cd",X"30", -- 1108
  X"28",X"7c",X"b5",X"ca",X"40",X"11",X"c1",X"e1", -- 1110
  X"e5",X"c5",X"e5",X"21",X"0b",X"00",X"39",X"cd", -- 1118
  X"d5",X"27",X"e5",X"3e",X"01",X"cd",X"22",X"1b", -- 1120
  X"c1",X"d1",X"cd",X"15",X"28",X"21",X"0d",X"00", -- 1128
  X"39",X"e5",X"cd",X"d5",X"27",X"11",X"02",X"00", -- 1130
  X"19",X"d1",X"cd",X"15",X"28",X"c3",X"84",X"11", -- 1138
  X"21",X"04",X"00",X"39",X"cd",X"c8",X"27",X"e5", -- 1140
  X"3e",X"01",X"cd",X"02",X"27",X"c1",X"cd",X"d5", -- 1148
  X"27",X"eb",X"21",X"02",X"00",X"cd",X"30",X"28", -- 1150
  X"7c",X"b5",X"ca",X"84",X"11",X"c1",X"e1",X"e5", -- 1158
  X"c5",X"e5",X"21",X"09",X"00",X"39",X"cd",X"d5", -- 1160
  X"27",X"e5",X"3e",X"01",X"cd",X"22",X"1b",X"c1", -- 1168
  X"d1",X"cd",X"15",X"28",X"21",X"0d",X"00",X"39", -- 1170
  X"e5",X"cd",X"d5",X"27",X"11",X"02",X"00",X"19", -- 1178
  X"d1",X"cd",X"15",X"28",X"21",X"0d",X"00",X"39", -- 1180
  X"cd",X"d5",X"27",X"33",X"c1",X"c1",X"c9",X"45", -- 1188
  X"52",X"52",X"4f",X"52",X"2d",X"00",X"21",X"5b", -- 1190
  X"00",X"e5",X"3e",X"01",X"cd",X"3e",X"1f",X"c1", -- 1198
  X"c1",X"e1",X"e5",X"c5",X"e5",X"3e",X"01",X"cd", -- 11a0
  X"6a",X"1c",X"c1",X"21",X"5d",X"00",X"e5",X"3e", -- 11a8
  X"01",X"cd",X"3e",X"1f",X"c1",X"c9",X"21",X"06", -- 11b0
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27", -- 11b8
  X"eb",X"21",X"00",X"00",X"cd",X"36",X"28",X"7c", -- 11c0
  X"b5",X"ca",X"0c",X"12",X"21",X"06",X"00",X"39", -- 11c8
  X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"e5",X"3e", -- 11d0
  X"01",X"cd",X"ef",X"14",X"c1",X"7c",X"b5",X"c2", -- 11d8
  X"fe",X"11",X"21",X"06",X"00",X"39",X"cd",X"d5", -- 11e0
  X"27",X"cd",X"c8",X"27",X"eb",X"21",X"2c",X"00", -- 11e8
  X"cd",X"30",X"28",X"7c",X"b5",X"c2",X"fe",X"11", -- 11f0
  X"21",X"00",X"00",X"c3",X"01",X"12",X"21",X"01", -- 11f8
  X"00",X"7c",X"b5",X"ca",X"0c",X"12",X"21",X"01", -- 1200
  X"00",X"c3",X"0f",X"12",X"21",X"00",X"00",X"7c", -- 1208
  X"b5",X"ca",X"25",X"12",X"21",X"06",X"00",X"39", -- 1210
  X"54",X"5d",X"cd",X"d5",X"27",X"23",X"cd",X"15", -- 1218
  X"28",X"2b",X"c3",X"b6",X"11",X"21",X"06",X"00", -- 1220
  X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"eb", -- 1228
  X"21",X"00",X"00",X"cd",X"36",X"28",X"7c",X"b5", -- 1230
  X"ca",X"70",X"12",X"21",X"06",X"00",X"39",X"cd", -- 1238
  X"d5",X"27",X"cd",X"c8",X"27",X"e5",X"3e",X"01", -- 1240
  X"cd",X"ef",X"14",X"c1",X"cd",X"9f",X"28",X"7c", -- 1248
  X"b5",X"ca",X"70",X"12",X"21",X"06",X"00",X"39", -- 1250
  X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"eb",X"21", -- 1258
  X"2c",X"00",X"cd",X"36",X"28",X"7c",X"b5",X"ca", -- 1260
  X"70",X"12",X"21",X"01",X"00",X"c3",X"73",X"12", -- 1268
  X"21",X"00",X"00",X"7c",X"b5",X"ca",X"9e",X"12", -- 1270
  X"21",X"04",X"00",X"39",X"54",X"5d",X"cd",X"d5", -- 1278
  X"27",X"23",X"cd",X"15",X"28",X"2b",X"e5",X"21", -- 1280
  X"08",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 1288
  X"23",X"cd",X"15",X"28",X"2b",X"cd",X"c8",X"27", -- 1290
  X"d1",X"7d",X"12",X"c3",X"25",X"12",X"21",X"04", -- 1298
  X"00",X"39",X"cd",X"d5",X"27",X"eb",X"21",X"00", -- 12a0
  X"00",X"7d",X"12",X"21",X"06",X"00",X"39",X"cd", -- 12a8
  X"d5",X"27",X"cd",X"c8",X"27",X"eb",X"21",X"00", -- 12b0
  X"00",X"cd",X"36",X"28",X"7c",X"b5",X"ca",X"dd", -- 12b8
  X"12",X"21",X"06",X"00",X"39",X"cd",X"d5",X"27", -- 12c0
  X"cd",X"c8",X"27",X"eb",X"21",X"20",X"00",X"cd", -- 12c8
  X"30",X"28",X"7c",X"b5",X"ca",X"dd",X"12",X"21", -- 12d0
  X"01",X"00",X"c3",X"e0",X"12",X"21",X"00",X"00", -- 12d8
  X"7c",X"b5",X"ca",X"f6",X"12",X"21",X"06",X"00", -- 12e0
  X"39",X"54",X"5d",X"cd",X"d5",X"27",X"23",X"cd", -- 12e8
  X"15",X"28",X"2b",X"c3",X"ab",X"12",X"21",X"06", -- 12f0
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27", -- 12f8
  X"7c",X"b5",X"ca",X"2b",X"13",X"21",X"02",X"00", -- 1300
  X"39",X"54",X"5d",X"cd",X"d5",X"27",X"23",X"cd", -- 1308
  X"15",X"28",X"2b",X"e5",X"21",X"08",X"00",X"39", -- 1310
  X"54",X"5d",X"cd",X"d5",X"27",X"23",X"cd",X"15", -- 1318
  X"28",X"2b",X"cd",X"c8",X"27",X"d1",X"7d",X"12", -- 1320
  X"c3",X"f6",X"12",X"c1",X"d1",X"d5",X"c5",X"21", -- 1328
  X"00",X"00",X"7d",X"12",X"c9",X"21",X"06",X"00", -- 1330
  X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"eb", -- 1338
  X"21",X"00",X"00",X"cd",X"36",X"28",X"7c",X"b5", -- 1340
  X"ca",X"67",X"13",X"21",X"06",X"00",X"39",X"cd", -- 1348
  X"d5",X"27",X"cd",X"c8",X"27",X"eb",X"21",X"20", -- 1350
  X"00",X"cd",X"30",X"28",X"7c",X"b5",X"ca",X"67", -- 1358
  X"13",X"21",X"01",X"00",X"c3",X"6a",X"13",X"21", -- 1360
  X"00",X"00",X"7c",X"b5",X"ca",X"80",X"13",X"21", -- 1368
  X"06",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 1370
  X"23",X"cd",X"15",X"28",X"2b",X"c3",X"35",X"13", -- 1378
  X"21",X"06",X"00",X"39",X"cd",X"d5",X"27",X"cd", -- 1380
  X"c8",X"27",X"eb",X"21",X"00",X"00",X"cd",X"36", -- 1388
  X"28",X"7c",X"b5",X"ca",X"b2",X"13",X"21",X"06", -- 1390
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27", -- 1398
  X"eb",X"21",X"2c",X"00",X"cd",X"36",X"28",X"7c", -- 13a0
  X"b5",X"ca",X"b2",X"13",X"21",X"01",X"00",X"c3", -- 13a8
  X"b5",X"13",X"21",X"00",X"00",X"7c",X"b5",X"ca", -- 13b0
  X"e0",X"13",X"21",X"04",X"00",X"39",X"54",X"5d", -- 13b8
  X"cd",X"d5",X"27",X"23",X"cd",X"15",X"28",X"2b", -- 13c0
  X"e5",X"21",X"08",X"00",X"39",X"54",X"5d",X"cd", -- 13c8
  X"d5",X"27",X"23",X"cd",X"15",X"28",X"2b",X"cd", -- 13d0
  X"c8",X"27",X"d1",X"7d",X"12",X"c3",X"80",X"13", -- 13d8
  X"21",X"04",X"00",X"39",X"cd",X"d5",X"27",X"eb", -- 13e0
  X"21",X"00",X"00",X"7d",X"12",X"21",X"06",X"00", -- 13e8
  X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"eb", -- 13f0
  X"21",X"00",X"00",X"cd",X"36",X"28",X"7c",X"b5", -- 13f8
  X"ca",X"1f",X"14",X"21",X"06",X"00",X"39",X"cd", -- 1400
  X"d5",X"27",X"cd",X"c8",X"27",X"eb",X"21",X"2c", -- 1408
  X"00",X"cd",X"30",X"28",X"7c",X"b5",X"ca",X"1f", -- 1410
  X"14",X"21",X"01",X"00",X"c3",X"22",X"14",X"21", -- 1418
  X"00",X"00",X"7c",X"b5",X"ca",X"35",X"14",X"21", -- 1420
  X"06",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 1428
  X"23",X"cd",X"15",X"28",X"2b",X"21",X"06",X"00", -- 1430
  X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"eb", -- 1438
  X"21",X"00",X"00",X"cd",X"36",X"28",X"7c",X"b5", -- 1440
  X"ca",X"67",X"14",X"21",X"06",X"00",X"39",X"cd", -- 1448
  X"d5",X"27",X"cd",X"c8",X"27",X"eb",X"21",X"20", -- 1450
  X"00",X"cd",X"30",X"28",X"7c",X"b5",X"ca",X"67", -- 1458
  X"14",X"21",X"01",X"00",X"c3",X"6a",X"14",X"21", -- 1460
  X"00",X"00",X"7c",X"b5",X"ca",X"80",X"14",X"21", -- 1468
  X"06",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 1470
  X"23",X"cd",X"15",X"28",X"2b",X"c3",X"35",X"14", -- 1478
  X"21",X"06",X"00",X"39",X"cd",X"d5",X"27",X"cd", -- 1480
  X"c8",X"27",X"7c",X"b5",X"ca",X"b5",X"14",X"21", -- 1488
  X"02",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 1490
  X"23",X"cd",X"15",X"28",X"2b",X"e5",X"21",X"08", -- 1498
  X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27",X"23", -- 14a0
  X"cd",X"15",X"28",X"2b",X"cd",X"c8",X"27",X"d1", -- 14a8
  X"7d",X"12",X"c3",X"80",X"14",X"c1",X"d1",X"d5", -- 14b0
  X"c5",X"21",X"00",X"00",X"7d",X"12",X"c9",X"21", -- 14b8
  X"02",X"00",X"39",X"cd",X"c8",X"27",X"eb",X"21", -- 14c0
  X"20",X"00",X"cd",X"4a",X"28",X"7c",X"b5",X"ca", -- 14c8
  X"eb",X"14",X"21",X"02",X"00",X"39",X"cd",X"c8", -- 14d0
  X"27",X"eb",X"21",X"7e",X"00",X"cd",X"43",X"28", -- 14d8
  X"7c",X"b5",X"ca",X"eb",X"14",X"21",X"01",X"00", -- 14e0
  X"c3",X"ee",X"14",X"21",X"00",X"00",X"c9",X"21", -- 14e8
  X"02",X"00",X"39",X"cd",X"c8",X"27",X"eb",X"21", -- 14f0
  X"20",X"00",X"cd",X"43",X"28",X"7c",X"b5",X"ca", -- 14f8
  X"5d",X"15",X"21",X"02",X"00",X"39",X"cd",X"c8", -- 1500
  X"27",X"eb",X"21",X"20",X"00",X"cd",X"30",X"28", -- 1508
  X"7c",X"b5",X"c2",X"4f",X"15",X"21",X"02",X"00", -- 1510
  X"39",X"cd",X"c8",X"27",X"eb",X"21",X"0d",X"00", -- 1518
  X"cd",X"43",X"28",X"7c",X"b5",X"ca",X"41",X"15", -- 1520
  X"21",X"02",X"00",X"39",X"cd",X"c8",X"27",X"eb", -- 1528
  X"21",X"09",X"00",X"cd",X"4a",X"28",X"7c",X"b5", -- 1530
  X"ca",X"41",X"15",X"21",X"01",X"00",X"c3",X"44", -- 1538
  X"15",X"21",X"00",X"00",X"7c",X"b5",X"c2",X"4f", -- 1540
  X"15",X"21",X"00",X"00",X"c3",X"52",X"15",X"21", -- 1548
  X"01",X"00",X"7c",X"b5",X"ca",X"5d",X"15",X"21", -- 1550
  X"01",X"00",X"c3",X"60",X"15",X"21",X"00",X"00", -- 1558
  X"c9",X"21",X"02",X"00",X"39",X"cd",X"c8",X"27", -- 1560
  X"eb",X"21",X"66",X"00",X"cd",X"43",X"28",X"7c", -- 1568
  X"b5",X"ca",X"8d",X"15",X"21",X"02",X"00",X"39", -- 1570
  X"cd",X"c8",X"27",X"eb",X"21",X"61",X"00",X"cd", -- 1578
  X"4a",X"28",X"7c",X"b5",X"ca",X"8d",X"15",X"21", -- 1580
  X"01",X"00",X"c3",X"90",X"15",X"21",X"00",X"00", -- 1588
  X"7c",X"b5",X"c2",X"03",X"16",X"21",X"02",X"00", -- 1590
  X"39",X"cd",X"c8",X"27",X"eb",X"21",X"46",X"00", -- 1598
  X"cd",X"43",X"28",X"7c",X"b5",X"ca",X"c1",X"15", -- 15a0
  X"21",X"02",X"00",X"39",X"cd",X"c8",X"27",X"eb", -- 15a8
  X"21",X"41",X"00",X"cd",X"4a",X"28",X"7c",X"b5", -- 15b0
  X"ca",X"c1",X"15",X"21",X"01",X"00",X"c3",X"c4", -- 15b8
  X"15",X"21",X"00",X"00",X"7c",X"b5",X"c2",X"03", -- 15c0
  X"16",X"21",X"02",X"00",X"39",X"cd",X"c8",X"27", -- 15c8
  X"eb",X"21",X"39",X"00",X"cd",X"43",X"28",X"7c", -- 15d0
  X"b5",X"ca",X"f5",X"15",X"21",X"02",X"00",X"39", -- 15d8
  X"cd",X"c8",X"27",X"eb",X"21",X"30",X"00",X"cd", -- 15e0
  X"4a",X"28",X"7c",X"b5",X"ca",X"f5",X"15",X"21", -- 15e8
  X"01",X"00",X"c3",X"f8",X"15",X"21",X"00",X"00", -- 15f0
  X"7c",X"b5",X"c2",X"03",X"16",X"21",X"00",X"00", -- 15f8
  X"c3",X"06",X"16",X"21",X"01",X"00",X"c9",X"c1", -- 1600
  X"e1",X"e5",X"c5",X"cd",X"c8",X"27",X"eb",X"21", -- 1608
  X"00",X"00",X"cd",X"30",X"28",X"7c",X"b5",X"c2", -- 1610
  X"3c",X"16",X"c1",X"e1",X"e5",X"c5",X"e5",X"21", -- 1618
  X"15",X"17",X"e5",X"3e",X"02",X"cd",X"54",X"17", -- 1620
  X"c1",X"c1",X"eb",X"21",X"00",X"00",X"cd",X"30", -- 1628
  X"28",X"7c",X"b5",X"c2",X"3c",X"16",X"21",X"00", -- 1630
  X"00",X"c3",X"3f",X"16",X"21",X"01",X"00",X"7c", -- 1638
  X"b5",X"ca",X"48",X"16",X"21",X"00",X"00",X"c9", -- 1640
  X"c1",X"e1",X"e5",X"c5",X"e5",X"21",X"19",X"17", -- 1648
  X"e5",X"3e",X"02",X"cd",X"54",X"17",X"c1",X"c1", -- 1650
  X"eb",X"21",X"00",X"00",X"cd",X"30",X"28",X"7c", -- 1658
  X"b5",X"c2",X"86",X"16",X"c1",X"e1",X"e5",X"c5", -- 1660
  X"e5",X"21",X"1d",X"17",X"e5",X"3e",X"02",X"cd", -- 1668
  X"54",X"17",X"c1",X"c1",X"eb",X"21",X"00",X"00", -- 1670
  X"cd",X"30",X"28",X"7c",X"b5",X"c2",X"86",X"16", -- 1678
  X"21",X"00",X"00",X"c3",X"89",X"16",X"21",X"01", -- 1680
  X"00",X"7c",X"b5",X"ca",X"92",X"16",X"21",X"00", -- 1688
  X"00",X"c9",X"c1",X"e1",X"e5",X"c5",X"e5",X"21", -- 1690
  X"20",X"17",X"e5",X"3e",X"02",X"cd",X"54",X"17", -- 1698
  X"c1",X"c1",X"eb",X"21",X"00",X"00",X"cd",X"30", -- 16a0
  X"28",X"7c",X"b5",X"c2",X"d0",X"16",X"c1",X"e1", -- 16a8
  X"e5",X"c5",X"e5",X"21",X"24",X"17",X"e5",X"3e", -- 16b0
  X"02",X"cd",X"54",X"17",X"c1",X"c1",X"eb",X"21", -- 16b8
  X"00",X"00",X"cd",X"30",X"28",X"7c",X"b5",X"c2", -- 16c0
  X"d0",X"16",X"21",X"00",X"00",X"c3",X"d3",X"16", -- 16c8
  X"21",X"01",X"00",X"7c",X"b5",X"ca",X"dc",X"16", -- 16d0
  X"21",X"00",X"00",X"c9",X"c1",X"e1",X"e5",X"c5", -- 16d8
  X"cd",X"c8",X"27",X"e5",X"3e",X"01",X"cd",X"61", -- 16e0
  X"15",X"c1",X"7c",X"b5",X"ca",X"00",X"17",X"21", -- 16e8
  X"02",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 16f0
  X"23",X"cd",X"15",X"28",X"2b",X"c3",X"dc",X"16", -- 16f8
  X"c1",X"e1",X"e5",X"c5",X"cd",X"c8",X"27",X"7c", -- 1700
  X"b5",X"c2",X"10",X"17",X"21",X"01",X"00",X"c9", -- 1708
  X"21",X"00",X"00",X"c9",X"c9",X"41",X"44",X"43", -- 1710
  X"00",X"41",X"44",X"44",X"00",X"43",X"43",X"00", -- 1718
  X"44",X"41",X"41",X"00",X"44",X"41",X"44",X"00", -- 1720
  X"21",X"04",X"00",X"39",X"54",X"5d",X"cd",X"d5", -- 1728
  X"27",X"23",X"cd",X"15",X"28",X"2b",X"e5",X"21", -- 1730
  X"04",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 1738
  X"23",X"cd",X"15",X"28",X"2b",X"cd",X"c8",X"27", -- 1740
  X"d1",X"7d",X"12",X"7c",X"b5",X"ca",X"53",X"17", -- 1748
  X"c3",X"28",X"17",X"c9",X"21",X"04",X"00",X"39", -- 1750
  X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"eb",X"c1", -- 1758
  X"e1",X"e5",X"c5",X"cd",X"c8",X"27",X"cd",X"30", -- 1760
  X"28",X"7c",X"b5",X"ca",X"9e",X"17",X"21",X"04", -- 1768
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27", -- 1770
  X"7c",X"b5",X"c2",X"81",X"17",X"21",X"00",X"00", -- 1778
  X"c9",X"21",X"04",X"00",X"39",X"54",X"5d",X"cd", -- 1780
  X"d5",X"27",X"23",X"cd",X"15",X"28",X"21",X"02", -- 1788
  X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27",X"23", -- 1790
  X"cd",X"15",X"28",X"c3",X"54",X"17",X"21",X"04", -- 1798
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27", -- 17a0
  X"eb",X"c1",X"e1",X"e5",X"c5",X"cd",X"c8",X"27", -- 17a8
  X"cd",X"8c",X"28",X"c9",X"21",X"f3",X"ff",X"39", -- 17b0
  X"f9",X"21",X"0b",X"00",X"39",X"eb",X"21",X"00", -- 17b8
  X"00",X"cd",X"15",X"28",X"21",X"0b",X"00",X"39", -- 17c0
  X"cd",X"d5",X"27",X"eb",X"21",X"08",X"00",X"cd", -- 17c8
  X"50",X"28",X"7c",X"b5",X"ca",X"01",X"18",X"c3", -- 17d0
  X"eb",X"17",X"21",X"0b",X"00",X"39",X"54",X"5d", -- 17d8
  X"cd",X"d5",X"27",X"23",X"cd",X"15",X"28",X"2b", -- 17e0
  X"c3",X"c4",X"17",X"21",X"00",X"00",X"39",X"eb", -- 17e8
  X"21",X"0b",X"00",X"39",X"cd",X"d5",X"27",X"19", -- 17f0
  X"eb",X"21",X"20",X"00",X"7d",X"12",X"c3",X"da", -- 17f8
  X"17",X"21",X"08",X"00",X"39",X"e5",X"21",X"13", -- 1800
  X"00",X"39",X"cd",X"d5",X"27",X"eb",X"21",X"00", -- 1808
  X"00",X"cd",X"4a",X"28",X"7c",X"b5",X"ca",X"1f", -- 1810
  X"18",X"21",X"2b",X"00",X"c3",X"22",X"18",X"21", -- 1818
  X"2d",X"00",X"d1",X"7d",X"12",X"21",X"0b",X"00", -- 1820
  X"39",X"eb",X"21",X"07",X"00",X"cd",X"15",X"28", -- 1828
  X"21",X"00",X"00",X"39",X"eb",X"21",X"0b",X"00", -- 1830
  X"39",X"cd",X"d5",X"27",X"19",X"e5",X"21",X"13", -- 1838
  X"00",X"39",X"cd",X"d5",X"27",X"eb",X"21",X"0a", -- 1840
  X"00",X"cd",X"33",X"27",X"eb",X"11",X"30",X"00", -- 1848
  X"19",X"d1",X"7d",X"12",X"21",X"11",X"00",X"39", -- 1850
  X"e5",X"21",X"13",X"00",X"39",X"cd",X"d5",X"27", -- 1858
  X"eb",X"21",X"0a",X"00",X"cd",X"33",X"27",X"d1", -- 1860
  X"cd",X"15",X"28",X"21",X"0b",X"00",X"39",X"54", -- 1868
  X"5d",X"cd",X"d5",X"27",X"2b",X"cd",X"15",X"28", -- 1870
  X"23",X"21",X"11",X"00",X"39",X"cd",X"d5",X"27", -- 1878
  X"af",X"b4",X"fa",X"8c",X"18",X"b5",X"ca",X"8c", -- 1880
  X"18",X"c3",X"30",X"18",X"21",X"00",X"00",X"39", -- 1888
  X"eb",X"21",X"0b",X"00",X"39",X"cd",X"d5",X"27", -- 1890
  X"19",X"eb",X"21",X"08",X"00",X"39",X"cd",X"c8", -- 1898
  X"27",X"7d",X"12",X"21",X"09",X"00",X"39",X"eb", -- 18a0
  X"21",X"00",X"00",X"cd",X"15",X"28",X"21",X"0b", -- 18a8
  X"00",X"39",X"cd",X"d5",X"27",X"eb",X"21",X"08", -- 18b0
  X"00",X"cd",X"50",X"28",X"7c",X"b5",X"ca",X"f8", -- 18b8
  X"18",X"21",X"0f",X"00",X"39",X"cd",X"d5",X"27", -- 18c0
  X"e5",X"21",X"0b",X"00",X"39",X"54",X"5d",X"cd", -- 18c8
  X"d5",X"27",X"23",X"cd",X"15",X"28",X"2b",X"d1", -- 18d0
  X"19",X"e5",X"21",X"02",X"00",X"39",X"e5",X"21", -- 18d8
  X"0f",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 18e0
  X"23",X"cd",X"15",X"28",X"2b",X"d1",X"19",X"cd", -- 18e8
  X"c8",X"27",X"d1",X"7d",X"12",X"c3",X"ae",X"18", -- 18f0
  X"21",X"0f",X"00",X"39",X"cd",X"d5",X"27",X"eb", -- 18f8
  X"21",X"09",X"00",X"39",X"cd",X"d5",X"27",X"19", -- 1900
  X"eb",X"21",X"00",X"00",X"7d",X"12",X"21",X"0d", -- 1908
  X"00",X"39",X"f9",X"c9",X"c5",X"c5",X"21",X"00", -- 1910
  X"00",X"39",X"e5",X"21",X"04",X"00",X"39",X"eb", -- 1918
  X"21",X"00",X"00",X"cd",X"15",X"28",X"d1",X"cd", -- 1920
  X"15",X"28",X"21",X"06",X"00",X"39",X"cd",X"d5", -- 1928
  X"27",X"cd",X"c8",X"27",X"eb",X"21",X"2b",X"00", -- 1930
  X"cd",X"30",X"28",X"7c",X"b5",X"c2",X"5c",X"19", -- 1938
  X"21",X"06",X"00",X"39",X"cd",X"d5",X"27",X"cd", -- 1940
  X"c8",X"27",X"eb",X"21",X"2d",X"00",X"cd",X"30", -- 1948
  X"28",X"7c",X"b5",X"c2",X"5c",X"19",X"21",X"00", -- 1950
  X"00",X"c3",X"5f",X"19",X"21",X"01",X"00",X"7c", -- 1958
  X"b5",X"ca",X"8e",X"19",X"21",X"06",X"00",X"39", -- 1960
  X"54",X"5d",X"cd",X"d5",X"27",X"23",X"cd",X"15", -- 1968
  X"28",X"2b",X"cd",X"c8",X"27",X"eb",X"21",X"2d", -- 1970
  X"00",X"cd",X"30",X"28",X"7c",X"b5",X"ca",X"8e", -- 1978
  X"19",X"21",X"00",X"00",X"39",X"eb",X"e1",X"e5", -- 1980
  X"cd",X"93",X"28",X"cd",X"15",X"28",X"21",X"06", -- 1988
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27", -- 1990
  X"7c",X"b5",X"ca",X"d1",X"19",X"21",X"02",X"00", -- 1998
  X"39",X"e5",X"21",X"04",X"00",X"39",X"cd",X"d5", -- 19a0
  X"27",X"11",X"0a",X"00",X"cd",X"13",X"27",X"e5", -- 19a8
  X"21",X"0a",X"00",X"39",X"54",X"5d",X"cd",X"d5", -- 19b0
  X"27",X"23",X"cd",X"15",X"28",X"2b",X"cd",X"c8", -- 19b8
  X"27",X"d1",X"19",X"eb",X"21",X"30",X"00",X"cd", -- 19c0
  X"8c",X"28",X"d1",X"cd",X"15",X"28",X"c3",X"8e", -- 19c8
  X"19",X"e1",X"e5",X"7c",X"b5",X"ca",X"e2",X"19", -- 19d0
  X"c1",X"e1",X"e5",X"c5",X"cd",X"93",X"28",X"c1", -- 19d8
  X"c1",X"c9",X"c1",X"e1",X"e5",X"c5",X"c1",X"c1", -- 19e0
  X"c9",X"c5",X"21",X"01",X"00",X"39",X"eb",X"21", -- 19e8
  X"00",X"00",X"7d",X"12",X"21",X"04",X"00",X"39", -- 19f0
  X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"7c",X"b5", -- 19f8
  X"ca",X"19",X"1b",X"21",X"04",X"00",X"39",X"cd", -- 1a00
  X"d5",X"27",X"cd",X"c8",X"27",X"eb",X"21",X"30", -- 1a08
  X"00",X"cd",X"4a",X"28",X"7c",X"b5",X"ca",X"35", -- 1a10
  X"1a",X"21",X"04",X"00",X"39",X"cd",X"d5",X"27", -- 1a18
  X"cd",X"c8",X"27",X"eb",X"21",X"39",X"00",X"cd", -- 1a20
  X"43",X"28",X"7c",X"b5",X"ca",X"35",X"1a",X"21", -- 1a28
  X"01",X"00",X"c3",X"38",X"1a",X"21",X"00",X"00", -- 1a30
  X"7c",X"b5",X"ca",X"4a",X"1a",X"21",X"00",X"00", -- 1a38
  X"39",X"eb",X"21",X"30",X"00",X"7d",X"12",X"c3", -- 1a40
  X"db",X"1a",X"21",X"04",X"00",X"39",X"cd",X"d5", -- 1a48
  X"27",X"cd",X"c8",X"27",X"eb",X"21",X"41",X"00", -- 1a50
  X"cd",X"4a",X"28",X"7c",X"b5",X"ca",X"7c",X"1a", -- 1a58
  X"21",X"04",X"00",X"39",X"cd",X"d5",X"27",X"cd", -- 1a60
  X"c8",X"27",X"eb",X"21",X"46",X"00",X"cd",X"43", -- 1a68
  X"28",X"7c",X"b5",X"ca",X"7c",X"1a",X"21",X"01", -- 1a70
  X"00",X"c3",X"7f",X"1a",X"21",X"00",X"00",X"7c", -- 1a78
  X"b5",X"ca",X"91",X"1a",X"21",X"00",X"00",X"39", -- 1a80
  X"eb",X"21",X"37",X"00",X"7d",X"12",X"c3",X"db", -- 1a88
  X"1a",X"21",X"04",X"00",X"39",X"cd",X"d5",X"27", -- 1a90
  X"cd",X"c8",X"27",X"eb",X"21",X"61",X"00",X"cd", -- 1a98
  X"4a",X"28",X"7c",X"b5",X"ca",X"c3",X"1a",X"21", -- 1aa0
  X"04",X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8", -- 1aa8
  X"27",X"eb",X"21",X"66",X"00",X"cd",X"43",X"28", -- 1ab0
  X"7c",X"b5",X"ca",X"c3",X"1a",X"21",X"01",X"00", -- 1ab8
  X"c3",X"c6",X"1a",X"21",X"00",X"00",X"7c",X"b5", -- 1ac0
  X"ca",X"d8",X"1a",X"21",X"00",X"00",X"39",X"eb", -- 1ac8
  X"21",X"57",X"00",X"7d",X"12",X"c3",X"db",X"1a", -- 1ad0
  X"c3",X"19",X"1b",X"21",X"01",X"00",X"39",X"e5", -- 1ad8
  X"21",X"03",X"00",X"39",X"cd",X"c8",X"27",X"eb", -- 1ae0
  X"21",X"04",X"00",X"cd",X"b9",X"27",X"eb",X"21", -- 1ae8
  X"06",X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8", -- 1af0
  X"27",X"19",X"eb",X"21",X"02",X"00",X"39",X"cd", -- 1af8
  X"c8",X"27",X"cd",X"8c",X"28",X"d1",X"7d",X"12", -- 1b00
  X"21",X"04",X"00",X"39",X"54",X"5d",X"cd",X"d5", -- 1b08
  X"27",X"23",X"cd",X"15",X"28",X"2b",X"c3",X"f4", -- 1b10
  X"19",X"21",X"01",X"00",X"39",X"cd",X"c8",X"27", -- 1b18
  X"c1",X"c9",X"c5",X"c5",X"21",X"02",X"00",X"39", -- 1b20
  X"eb",X"21",X"00",X"00",X"cd",X"15",X"28",X"21", -- 1b28
  X"06",X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8", -- 1b30
  X"27",X"7c",X"b5",X"ca",X"55",X"1c",X"21",X"06", -- 1b38
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27", -- 1b40
  X"eb",X"21",X"30",X"00",X"cd",X"4a",X"28",X"7c", -- 1b48
  X"b5",X"ca",X"70",X"1b",X"21",X"06",X"00",X"39", -- 1b50
  X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"eb",X"21", -- 1b58
  X"39",X"00",X"cd",X"43",X"28",X"7c",X"b5",X"ca", -- 1b60
  X"70",X"1b",X"21",X"01",X"00",X"c3",X"73",X"1b", -- 1b68
  X"21",X"00",X"00",X"7c",X"b5",X"ca",X"86",X"1b", -- 1b70
  X"21",X"00",X"00",X"39",X"eb",X"21",X"30",X"00", -- 1b78
  X"cd",X"15",X"28",X"c3",X"19",X"1c",X"21",X"06", -- 1b80
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27", -- 1b88
  X"eb",X"21",X"41",X"00",X"cd",X"4a",X"28",X"7c", -- 1b90
  X"b5",X"ca",X"b8",X"1b",X"21",X"06",X"00",X"39", -- 1b98
  X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"eb",X"21", -- 1ba0
  X"46",X"00",X"cd",X"43",X"28",X"7c",X"b5",X"ca", -- 1ba8
  X"b8",X"1b",X"21",X"01",X"00",X"c3",X"bb",X"1b", -- 1bb0
  X"21",X"00",X"00",X"7c",X"b5",X"ca",X"ce",X"1b", -- 1bb8
  X"21",X"00",X"00",X"39",X"eb",X"21",X"37",X"00", -- 1bc0
  X"cd",X"15",X"28",X"c3",X"19",X"1c",X"21",X"06", -- 1bc8
  X"00",X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27", -- 1bd0
  X"eb",X"21",X"61",X"00",X"cd",X"4a",X"28",X"7c", -- 1bd8
  X"b5",X"ca",X"00",X"1c",X"21",X"06",X"00",X"39", -- 1be0
  X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"eb",X"21", -- 1be8
  X"66",X"00",X"cd",X"43",X"28",X"7c",X"b5",X"ca", -- 1bf0
  X"00",X"1c",X"21",X"01",X"00",X"c3",X"03",X"1c", -- 1bf8
  X"21",X"00",X"00",X"7c",X"b5",X"ca",X"16",X"1c", -- 1c00
  X"21",X"00",X"00",X"39",X"eb",X"21",X"57",X"00", -- 1c08
  X"cd",X"15",X"28",X"c3",X"19",X"1c",X"c3",X"55", -- 1c10
  X"1c",X"21",X"02",X"00",X"39",X"e5",X"21",X"04", -- 1c18
  X"00",X"39",X"cd",X"d5",X"27",X"eb",X"21",X"04", -- 1c20
  X"00",X"cd",X"b9",X"27",X"eb",X"21",X"08",X"00", -- 1c28
  X"39",X"cd",X"d5",X"27",X"cd",X"c8",X"27",X"19", -- 1c30
  X"eb",X"c1",X"e1",X"e5",X"c5",X"cd",X"8c",X"28", -- 1c38
  X"d1",X"cd",X"15",X"28",X"21",X"06",X"00",X"39", -- 1c40
  X"54",X"5d",X"cd",X"d5",X"27",X"23",X"cd",X"15", -- 1c48
  X"28",X"2b",X"c3",X"2f",X"1b",X"c1",X"e1",X"e5", -- 1c50
  X"c5",X"c1",X"c1",X"c9",X"21",X"67",X"1c",X"e5", -- 1c58
  X"3e",X"01",X"cd",X"ef",X"1d",X"c1",X"c9",X"0d", -- 1c60
  X"0a",X"00",X"21",X"f8",X"ff",X"39",X"f9",X"21", -- 1c68
  X"00",X"00",X"39",X"eb",X"21",X"03",X"00",X"cd", -- 1c70
  X"15",X"28",X"e1",X"e5",X"af",X"b4",X"fa",X"10", -- 1c78
  X"1d",X"c3",X"95",X"1c",X"21",X"00",X"00",X"39", -- 1c80
  X"54",X"5d",X"cd",X"d5",X"27",X"2b",X"cd",X"15", -- 1c88
  X"28",X"23",X"c3",X"7a",X"1c",X"21",X"07",X"00", -- 1c90
  X"39",X"e5",X"21",X"0c",X"00",X"39",X"cd",X"d5", -- 1c98
  X"27",X"eb",X"21",X"0f",X"00",X"cd",X"29",X"28", -- 1ca0
  X"d1",X"7d",X"12",X"21",X"0a",X"00",X"39",X"e5", -- 1ca8
  X"21",X"0c",X"00",X"39",X"cd",X"d5",X"27",X"eb", -- 1cb0
  X"21",X"04",X"00",X"cd",X"ab",X"27",X"eb",X"21", -- 1cb8
  X"ff",X"0f",X"cd",X"29",X"28",X"d1",X"cd",X"15", -- 1cc0
  X"28",X"21",X"07",X"00",X"39",X"cd",X"c8",X"27", -- 1cc8
  X"eb",X"21",X"0a",X"00",X"cd",X"50",X"28",X"7c", -- 1cd0
  X"b5",X"ca",X"f6",X"1c",X"21",X"02",X"00",X"39", -- 1cd8
  X"eb",X"e1",X"e5",X"19",X"e5",X"21",X"09",X"00", -- 1ce0
  X"39",X"cd",X"c8",X"27",X"11",X"30",X"00",X"19", -- 1ce8
  X"d1",X"7d",X"12",X"c3",X"0d",X"1d",X"21",X"02", -- 1cf0
  X"00",X"39",X"eb",X"e1",X"e5",X"19",X"e5",X"21", -- 1cf8
  X"09",X"00",X"39",X"cd",X"c8",X"27",X"11",X"37", -- 1d00
  X"00",X"19",X"d1",X"7d",X"12",X"c3",X"84",X"1c", -- 1d08
  X"21",X"02",X"00",X"39",X"11",X"04",X"00",X"19", -- 1d10
  X"eb",X"21",X"00",X"00",X"7d",X"12",X"21",X"02", -- 1d18
  X"00",X"39",X"e5",X"3e",X"01",X"cd",X"ef",X"1d", -- 1d20
  X"c1",X"21",X"08",X"00",X"39",X"f9",X"c9",X"c5", -- 1d28
  X"c5",X"c5",X"21",X"00",X"00",X"39",X"eb",X"21", -- 1d30
  X"01",X"00",X"cd",X"15",X"28",X"e1",X"e5",X"af", -- 1d38
  X"b4",X"fa",X"d2",X"1d",X"c3",X"58",X"1d",X"21", -- 1d40
  X"00",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 1d48
  X"2b",X"cd",X"15",X"28",X"23",X"c3",X"3d",X"1d", -- 1d50
  X"21",X"05",X"00",X"39",X"e5",X"21",X"0a",X"00", -- 1d58
  X"39",X"cd",X"c8",X"27",X"eb",X"21",X"0f",X"00", -- 1d60
  X"cd",X"29",X"28",X"d1",X"7d",X"12",X"21",X"08", -- 1d68
  X"00",X"39",X"e5",X"21",X"0a",X"00",X"39",X"cd", -- 1d70
  X"c8",X"27",X"eb",X"21",X"04",X"00",X"cd",X"ab", -- 1d78
  X"27",X"eb",X"21",X"ff",X"0f",X"cd",X"29",X"28", -- 1d80
  X"d1",X"7d",X"12",X"21",X"05",X"00",X"39",X"cd", -- 1d88
  X"c8",X"27",X"eb",X"21",X"0a",X"00",X"cd",X"50", -- 1d90
  X"28",X"7c",X"b5",X"ca",X"b8",X"1d",X"21",X"02", -- 1d98
  X"00",X"39",X"eb",X"e1",X"e5",X"19",X"e5",X"21", -- 1da0
  X"07",X"00",X"39",X"cd",X"c8",X"27",X"11",X"30", -- 1da8
  X"00",X"19",X"d1",X"7d",X"12",X"c3",X"cf",X"1d", -- 1db0
  X"21",X"02",X"00",X"39",X"eb",X"e1",X"e5",X"19", -- 1db8
  X"e5",X"21",X"07",X"00",X"39",X"cd",X"c8",X"27", -- 1dc0
  X"11",X"37",X"00",X"19",X"d1",X"7d",X"12",X"c3", -- 1dc8
  X"47",X"1d",X"21",X"02",X"00",X"39",X"11",X"02", -- 1dd0
  X"00",X"19",X"eb",X"21",X"00",X"00",X"7d",X"12", -- 1dd8
  X"21",X"02",X"00",X"39",X"e5",X"3e",X"01",X"cd", -- 1de0
  X"ef",X"1d",X"c1",X"c1",X"c1",X"c1",X"c9",X"c1", -- 1de8
  X"e1",X"e5",X"c5",X"cd",X"c8",X"27",X"7c",X"b5", -- 1df0
  X"ca",X"16",X"1e",X"21",X"02",X"00",X"39",X"54", -- 1df8
  X"5d",X"cd",X"d5",X"27",X"23",X"cd",X"15",X"28", -- 1e00
  X"2b",X"cd",X"c8",X"27",X"e5",X"3e",X"01",X"cd", -- 1e08
  X"3e",X"1f",X"c1",X"c3",X"ef",X"1d",X"c9",X"3b", -- 1e10
  X"c5",X"21",X"00",X"00",X"39",X"eb",X"21",X"00", -- 1e18
  X"00",X"cd",X"15",X"28",X"21",X"02",X"00",X"39", -- 1e20
  X"e5",X"af",X"cd",X"48",X"1f",X"d1",X"7d",X"12", -- 1e28
  X"eb",X"21",X"0d",X"00",X"cd",X"36",X"28",X"7c", -- 1e30
  X"b5",X"ca",X"1b",X"1f",X"21",X"02",X"00",X"39", -- 1e38
  X"cd",X"c8",X"27",X"eb",X"21",X"09",X"00",X"cd", -- 1e40
  X"30",X"28",X"7c",X"b5",X"ca",X"59",X"1e",X"21", -- 1e48
  X"02",X"00",X"39",X"eb",X"21",X"20",X"00",X"7d", -- 1e50
  X"12",X"21",X"02",X"00",X"39",X"cd",X"c8",X"27", -- 1e58
  X"eb",X"21",X"08",X"00",X"cd",X"30",X"28",X"7c", -- 1e60
  X"b5",X"ca",X"7f",X"1e",X"d1",X"d5",X"21",X"00", -- 1e68
  X"00",X"cd",X"3c",X"28",X"7c",X"b5",X"ca",X"7f", -- 1e70
  X"1e",X"21",X"01",X"00",X"c3",X"82",X"1e",X"21", -- 1e78
  X"00",X"00",X"7c",X"b5",X"ca",X"b6",X"1e",X"21", -- 1e80
  X"00",X"00",X"39",X"54",X"5d",X"cd",X"d5",X"27", -- 1e88
  X"2b",X"cd",X"15",X"28",X"23",X"21",X"08",X"00", -- 1e90
  X"e5",X"3e",X"01",X"cd",X"3e",X"1f",X"c1",X"21", -- 1e98
  X"20",X"00",X"e5",X"3e",X"01",X"cd",X"3e",X"1f", -- 1ea0
  X"c1",X"21",X"08",X"00",X"e5",X"3e",X"01",X"cd", -- 1ea8
  X"3e",X"1f",X"c1",X"c3",X"18",X"1f",X"21",X"02", -- 1eb0
  X"00",X"39",X"cd",X"c8",X"27",X"e5",X"3e",X"01", -- 1eb8
  X"cd",X"bf",X"14",X"c1",X"7c",X"b5",X"ca",X"e0", -- 1ec0
  X"1e",X"d1",X"d5",X"21",X"05",X"00",X"39",X"cd", -- 1ec8
  X"d5",X"27",X"cd",X"50",X"28",X"7c",X"b5",X"ca", -- 1ed0
  X"e0",X"1e",X"21",X"01",X"00",X"c3",X"e3",X"1e", -- 1ed8
  X"21",X"00",X"00",X"7c",X"b5",X"ca",X"18",X"1f", -- 1ee0
  X"21",X"07",X"00",X"39",X"cd",X"d5",X"27",X"e5", -- 1ee8
  X"21",X"02",X"00",X"39",X"54",X"5d",X"cd",X"d5", -- 1ef0
  X"27",X"23",X"cd",X"15",X"28",X"2b",X"d1",X"19", -- 1ef8
  X"eb",X"21",X"02",X"00",X"39",X"cd",X"c8",X"27", -- 1f00
  X"7d",X"12",X"21",X"02",X"00",X"39",X"cd",X"c8", -- 1f08
  X"27",X"e5",X"3e",X"01",X"cd",X"3e",X"1f",X"c1", -- 1f10
  X"c3",X"24",X"1e",X"21",X"07",X"00",X"39",X"cd", -- 1f18
  X"d5",X"27",X"eb",X"e1",X"e5",X"19",X"eb",X"21", -- 1f20
  X"00",X"00",X"7d",X"12",X"af",X"cd",X"5c",X"1c", -- 1f28
  X"33",X"c1",X"c9",X"c1",X"d1",X"d5",X"c5",X"21", -- 1f30
  X"3d",X"1f",X"e5",X"eb",X"e9",X"c9",X"c1",X"d1", -- 1f38
  X"d5",X"c5",X"0e",X"02",X"cd",X"05",X"00",X"c9", -- 1f40
  X"0e",X"06",X"1e",X"ff",X"cd",X"05",X"00",X"fe", -- 1f48
  X"00",X"ca",X"48",X"1f",X"fe",X"61",X"da",X"60", -- 1f50
  X"1f",X"fe",X"7b",X"d2",X"60",X"1f",X"e6",X"df", -- 1f58
  X"26",X"00",X"6f",X"c9",X"0e",X"00",X"cd",X"05", -- 1f60
  X"00",X"c9",X"3f",X"00",X"41",X"43",X"49",X"00", -- 1f68
  X"41",X"44",X"43",X"00",X"41",X"44",X"44",X"00", -- 1f70
  X"41",X"44",X"49",X"00",X"41",X"4e",X"41",X"00", -- 1f78
  X"41",X"4e",X"49",X"00",X"43",X"41",X"4c",X"4c", -- 1f80
  X"00",X"43",X"43",X"00",X"43",X"4d",X"00",X"43", -- 1f88
  X"4d",X"41",X"00",X"43",X"4d",X"43",X"00",X"43", -- 1f90
  X"4d",X"50",X"00",X"43",X"4e",X"5a",X"00",X"43", -- 1f98
  X"50",X"00",X"43",X"50",X"45",X"00",X"43",X"50", -- 1fa0
  X"49",X"00",X"43",X"50",X"4f",X"00",X"43",X"5a", -- 1fa8
  X"00",X"44",X"41",X"41",X"00",X"44",X"41",X"44", -- 1fb0
  X"00",X"44",X"43",X"52",X"00",X"44",X"43",X"58", -- 1fb8
  X"00",X"44",X"49",X"00",X"45",X"49",X"00",X"48", -- 1fc0
  X"4c",X"54",X"00",X"49",X"4e",X"00",X"49",X"4e", -- 1fc8
  X"52",X"00",X"49",X"4e",X"58",X"00",X"4a",X"43", -- 1fd0
  X"00",X"4a",X"4e",X"43",X"00",X"4a",X"4d",X"00", -- 1fd8
  X"4a",X"4d",X"50",X"00",X"4a",X"4e",X"5a",X"00", -- 1fe0
  X"4a",X"50",X"00",X"4a",X"50",X"45",X"00",X"4a", -- 1fe8
  X"50",X"4f",X"00",X"4a",X"5a",X"00",X"4c",X"44", -- 1ff0
  X"41",X"00",X"4c",X"44",X"41",X"58",X"00",X"4c", -- 1ff8
  X"48",X"4c",X"44",X"00",X"4c",X"58",X"49",X"00", -- 2000
  X"4d",X"4f",X"56",X"00",X"4d",X"56",X"49",X"00", -- 2008
  X"4e",X"4f",X"50",X"00",X"4f",X"52",X"41",X"00", -- 2010
  X"4f",X"52",X"49",X"00",X"4f",X"55",X"54",X"00", -- 2018
  X"50",X"43",X"48",X"4c",X"00",X"50",X"4f",X"50", -- 2020
  X"00",X"50",X"55",X"53",X"48",X"00",X"52",X"41", -- 2028
  X"4c",X"00",X"52",X"41",X"52",X"00",X"52",X"43", -- 2030
  X"00",X"52",X"45",X"54",X"00",X"52",X"4c",X"43", -- 2038
  X"00",X"52",X"4d",X"00",X"52",X"4e",X"43",X"00", -- 2040
  X"52",X"4e",X"5a",X"00",X"52",X"50",X"00",X"52", -- 2048
  X"50",X"45",X"00",X"52",X"50",X"4f",X"00",X"52", -- 2050
  X"52",X"43",X"00",X"52",X"53",X"54",X"30",X"00", -- 2058
  X"52",X"53",X"54",X"31",X"00",X"52",X"53",X"54", -- 2060
  X"32",X"00",X"52",X"53",X"54",X"33",X"00",X"52", -- 2068
  X"53",X"54",X"34",X"00",X"52",X"53",X"54",X"35", -- 2070
  X"00",X"52",X"53",X"54",X"36",X"00",X"52",X"53", -- 2078
  X"54",X"37",X"00",X"52",X"5a",X"00",X"53",X"42", -- 2080
  X"42",X"00",X"53",X"42",X"49",X"00",X"53",X"48", -- 2088
  X"4c",X"44",X"00",X"53",X"50",X"48",X"4c",X"00", -- 2090
  X"53",X"54",X"41",X"00",X"53",X"54",X"41",X"58", -- 2098
  X"00",X"53",X"54",X"43",X"00",X"53",X"55",X"42", -- 20a0
  X"00",X"53",X"55",X"49",X"00",X"58",X"43",X"48", -- 20a8
  X"47",X"00",X"58",X"52",X"41",X"00",X"58",X"52", -- 20b0
  X"49",X"00",X"58",X"54",X"48",X"4c",X"00",X"43", -- 20b8
  X"4e",X"43",X"00",X"10",X"20",X"04",X"20",X"9c", -- 20c0
  X"20",X"d2",X"1f",X"ce",X"1f",X"b9",X"1f",X"0c", -- 20c8
  X"20",X"3d",X"20",X"6a",X"1f",X"b5",X"1f",X"fa", -- 20d0
  X"1f",X"bd",X"1f",X"ce",X"1f",X"b9",X"1f",X"0c", -- 20d8
  X"20",X"57",X"20",X"6a",X"1f",X"04",X"20",X"9c", -- 20e0
  X"20",X"d2",X"1f",X"ce",X"1f",X"b9",X"1f",X"0c", -- 20e8
  X"20",X"2e",X"20",X"6a",X"1f",X"b5",X"1f",X"fa", -- 20f0
  X"1f",X"bd",X"1f",X"ce",X"1f",X"b9",X"1f",X"0c", -- 20f8
  X"20",X"32",X"20",X"6a",X"1f",X"04",X"20",X"8e", -- 2100
  X"20",X"d2",X"1f",X"ce",X"1f",X"b9",X"1f",X"0c", -- 2108
  X"20",X"b1",X"1f",X"6a",X"1f",X"b5",X"1f",X"ff", -- 2110
  X"1f",X"bd",X"1f",X"ce",X"1f",X"b9",X"1f",X"0c", -- 2118
  X"20",X"8f",X"1f",X"6a",X"1f",X"04",X"20",X"98", -- 2120
  X"20",X"d2",X"1f",X"ce",X"1f",X"b9",X"1f",X"0c", -- 2128
  X"20",X"a1",X"20",X"6a",X"1f",X"b5",X"1f",X"f6", -- 2130
  X"1f",X"bd",X"1f",X"ce",X"1f",X"b9",X"1f",X"0c", -- 2138
  X"20",X"93",X"1f",X"08",X"20",X"08",X"20",X"08", -- 2140
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 2148
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 2150
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 2158
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 2160
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 2168
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 2170
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 2178
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 2180
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 2188
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 2190
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 2198
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 21a0
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"c7", -- 21a8
  X"1f",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 21b0
  X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"08", -- 21b8
  X"20",X"08",X"20",X"74",X"1f",X"74",X"1f",X"74", -- 21c0
  X"1f",X"74",X"1f",X"74",X"1f",X"74",X"1f",X"74", -- 21c8
  X"1f",X"74",X"1f",X"70",X"1f",X"70",X"1f",X"70", -- 21d0
  X"1f",X"70",X"1f",X"70",X"1f",X"70",X"1f",X"70", -- 21d8
  X"1f",X"70",X"1f",X"a5",X"20",X"a5",X"20",X"a5", -- 21e0
  X"20",X"a5",X"20",X"a5",X"20",X"a5",X"20",X"a5", -- 21e8
  X"20",X"a5",X"20",X"86",X"20",X"86",X"20",X"86", -- 21f0
  X"20",X"86",X"20",X"86",X"20",X"86",X"20",X"86", -- 21f8
  X"20",X"86",X"20",X"7c",X"1f",X"7c",X"1f",X"7c", -- 2200
  X"1f",X"7c",X"1f",X"7c",X"1f",X"7c",X"1f",X"7c", -- 2208
  X"1f",X"7c",X"1f",X"b2",X"20",X"b2",X"20",X"b2", -- 2210
  X"20",X"b2",X"20",X"b2",X"20",X"b2",X"20",X"b2", -- 2218
  X"20",X"b2",X"20",X"14",X"20",X"14",X"20",X"14", -- 2220
  X"20",X"14",X"20",X"14",X"20",X"14",X"20",X"14", -- 2228
  X"20",X"14",X"20",X"97",X"1f",X"97",X"1f",X"97", -- 2230
  X"1f",X"97",X"1f",X"97",X"1f",X"97",X"1f",X"97", -- 2238
  X"1f",X"97",X"1f",X"48",X"20",X"25",X"20",X"e4", -- 2240
  X"1f",X"e0",X"1f",X"9b",X"1f",X"29",X"20",X"78", -- 2248
  X"1f",X"5b",X"20",X"83",X"20",X"39",X"20",X"f3", -- 2250
  X"1f",X"6a",X"1f",X"ae",X"1f",X"84",X"1f",X"6c", -- 2258
  X"1f",X"60",X"20",X"44",X"20",X"25",X"20",X"d9", -- 2260
  X"1f",X"1c",X"20",X"bf",X"20",X"29",X"20",X"a9", -- 2268
  X"20",X"65",X"20",X"36",X"20",X"6a",X"1f",X"d6", -- 2270
  X"1f",X"cb",X"1f",X"89",X"1f",X"6a",X"1f",X"8a", -- 2278
  X"20",X"6a",X"20",X"53",X"20",X"25",X"20",X"ef", -- 2280
  X"1f",X"ba",X"20",X"aa",X"1f",X"29",X"20",X"80", -- 2288
  X"1f",X"6f",X"20",X"4f",X"20",X"20",X"20",X"eb", -- 2290
  X"1f",X"ad",X"20",X"a2",X"1f",X"6a",X"1f",X"b6", -- 2298
  X"20",X"74",X"20",X"4c",X"20",X"25",X"20",X"e8", -- 22a0
  X"1f",X"c1",X"1f",X"9f",X"1f",X"29",X"20",X"18", -- 22a8
  X"20",X"79",X"20",X"41",X"20",X"93",X"20",X"dd", -- 22b0
  X"1f",X"c4",X"1f",X"8c",X"1f",X"6a",X"1f",X"a6", -- 22b8
  X"1f",X"7e",X"20",X"00",X"00",X"01",X"00",X"02", -- 22c0
  X"00",X"42",X"00",X"43",X"00",X"44",X"00",X"45", -- 22c8
  X"00",X"48",X"00",X"4c",X"00",X"4d",X"00",X"41", -- 22d0
  X"00",X"50",X"53",X"57",X"00",X"53",X"50",X"00", -- 22d8
  X"c3",X"22",X"c9",X"22",X"c9",X"22",X"c9",X"22", -- 22e0
  X"c9",X"22",X"c9",X"22",X"c9",X"22",X"c3",X"22", -- 22e8
  X"c3",X"22",X"c9",X"22",X"c9",X"22",X"c9",X"22", -- 22f0
  X"cb",X"22",X"cb",X"22",X"cb",X"22",X"c3",X"22", -- 22f8
  X"c3",X"22",X"cd",X"22",X"cd",X"22",X"cd",X"22", -- 2300
  X"cd",X"22",X"cd",X"22",X"cd",X"22",X"c3",X"22", -- 2308
  X"c3",X"22",X"cd",X"22",X"cd",X"22",X"cd",X"22", -- 2310
  X"cf",X"22",X"cf",X"22",X"cf",X"22",X"c3",X"22", -- 2318
  X"c3",X"22",X"d1",X"22",X"c7",X"22",X"d1",X"22", -- 2320
  X"d1",X"22",X"d1",X"22",X"d1",X"22",X"c3",X"22", -- 2328
  X"c3",X"22",X"d1",X"22",X"c7",X"22",X"d1",X"22", -- 2330
  X"d3",X"22",X"d3",X"22",X"d3",X"22",X"c3",X"22", -- 2338
  X"c3",X"22",X"dd",X"22",X"c7",X"22",X"dd",X"22", -- 2340
  X"d5",X"22",X"d5",X"22",X"d5",X"22",X"c3",X"22", -- 2348
  X"c3",X"22",X"dd",X"22",X"c7",X"22",X"dd",X"22", -- 2350
  X"d7",X"22",X"d7",X"22",X"d7",X"22",X"c3",X"22", -- 2358
  X"c9",X"22",X"c9",X"22",X"c9",X"22",X"c9",X"22", -- 2360
  X"c9",X"22",X"c9",X"22",X"c9",X"22",X"c9",X"22", -- 2368
  X"cb",X"22",X"cb",X"22",X"cb",X"22",X"cb",X"22", -- 2370
  X"cb",X"22",X"cb",X"22",X"cb",X"22",X"cb",X"22", -- 2378
  X"cd",X"22",X"cd",X"22",X"cd",X"22",X"cd",X"22", -- 2380
  X"cd",X"22",X"cd",X"22",X"cd",X"22",X"cd",X"22", -- 2388
  X"cf",X"22",X"cf",X"22",X"cf",X"22",X"cf",X"22", -- 2390
  X"cf",X"22",X"cf",X"22",X"cf",X"22",X"cf",X"22", -- 2398
  X"d1",X"22",X"d1",X"22",X"d1",X"22",X"d1",X"22", -- 23a0
  X"d1",X"22",X"d1",X"22",X"d1",X"22",X"d1",X"22", -- 23a8
  X"d3",X"22",X"d3",X"22",X"d3",X"22",X"d3",X"22", -- 23b0
  X"d3",X"22",X"d3",X"22",X"d3",X"22",X"d3",X"22", -- 23b8
  X"d5",X"22",X"d5",X"22",X"d5",X"22",X"d5",X"22", -- 23c0
  X"d5",X"22",X"d5",X"22",X"c3",X"22",X"d5",X"22", -- 23c8
  X"d7",X"22",X"d7",X"22",X"d7",X"22",X"d7",X"22", -- 23d0
  X"d7",X"22",X"d7",X"22",X"d7",X"22",X"d7",X"22", -- 23d8
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 23e0
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 23e8
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 23f0
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 23f8
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 2400
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 2408
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 2410
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 2418
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 2420
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 2428
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 2430
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 2438
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 2440
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 2448
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 2450
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 2458
  X"c3",X"22",X"c9",X"22",X"c7",X"22",X"c7",X"22", -- 2460
  X"c7",X"22",X"c9",X"22",X"c5",X"22",X"c3",X"22", -- 2468
  X"c3",X"22",X"c3",X"22",X"c7",X"22",X"c7",X"22", -- 2470
  X"c7",X"22",X"c7",X"22",X"c5",X"22",X"c3",X"22", -- 2478
  X"c3",X"22",X"cd",X"22",X"c7",X"22",X"c5",X"22", -- 2480
  X"c7",X"22",X"cd",X"22",X"c5",X"22",X"c3",X"22", -- 2488
  X"c3",X"22",X"c3",X"22",X"c7",X"22",X"c5",X"22", -- 2490
  X"c7",X"22",X"c7",X"22",X"c5",X"22",X"c3",X"22", -- 2498
  X"c3",X"22",X"d1",X"22",X"c7",X"22",X"c3",X"22", -- 24a0
  X"c7",X"22",X"d1",X"22",X"c5",X"22",X"c3",X"22", -- 24a8
  X"c3",X"22",X"c3",X"22",X"c7",X"22",X"c3",X"22", -- 24b0
  X"c7",X"22",X"c7",X"22",X"c5",X"22",X"c3",X"22", -- 24b8
  X"c3",X"22",X"d9",X"22",X"c7",X"22",X"c3",X"22", -- 24c0
  X"c7",X"22",X"d9",X"22",X"c5",X"22",X"c3",X"22", -- 24c8
  X"c3",X"22",X"c3",X"22",X"c7",X"22",X"c3",X"22", -- 24d0
  X"c7",X"22",X"c7",X"22",X"c5",X"22",X"c3",X"22", -- 24d8
  X"c3",X"22",X"c7",X"22",X"c3",X"22",X"c3",X"22", -- 24e0
  X"c3",X"22",X"c3",X"22",X"c5",X"22",X"c3",X"22", -- 24e8
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 24f0
  X"c3",X"22",X"c3",X"22",X"c5",X"22",X"c3",X"22", -- 24f8
  X"c3",X"22",X"c7",X"22",X"c3",X"22",X"c3",X"22", -- 2500
  X"c3",X"22",X"c3",X"22",X"c5",X"22",X"c3",X"22", -- 2508
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2510
  X"c3",X"22",X"c3",X"22",X"c5",X"22",X"c3",X"22", -- 2518
  X"c3",X"22",X"c7",X"22",X"c3",X"22",X"c3",X"22", -- 2520
  X"c3",X"22",X"c3",X"22",X"c5",X"22",X"c3",X"22", -- 2528
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2530
  X"c3",X"22",X"c3",X"22",X"c5",X"22",X"c3",X"22", -- 2538
  X"c3",X"22",X"c7",X"22",X"c3",X"22",X"c3",X"22", -- 2540
  X"c3",X"22",X"c3",X"22",X"c5",X"22",X"c3",X"22", -- 2548
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2550
  X"c3",X"22",X"c3",X"22",X"c5",X"22",X"c3",X"22", -- 2558
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 2560
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 2568
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 2570
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 2578
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 2580
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 2588
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 2590
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 2598
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 25a0
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 25a8
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 25b0
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 25b8
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 25c0
  X"d1",X"22",X"d3",X"22",X"c3",X"22",X"d7",X"22", -- 25c8
  X"c9",X"22",X"cb",X"22",X"cd",X"22",X"cf",X"22", -- 25d0
  X"d1",X"22",X"d3",X"22",X"d5",X"22",X"d7",X"22", -- 25d8
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 25e0
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 25e8
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 25f0
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 25f8
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2600
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2608
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2610
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2618
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2620
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2628
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2630
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2638
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2640
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2648
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2650
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2658
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2660
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2668
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2670
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2678
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2680
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2688
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2690
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 2698
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 26a0
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 26a8
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 26b0
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 26b8
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 26c0
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 26c8
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 26d0
  X"c3",X"22",X"c3",X"22",X"c3",X"22",X"c3",X"22", -- 26d8
  X"d1",X"c1",X"c5",X"d5",X"11",X"c3",X"20",X"26", -- 26e0
  X"00",X"69",X"29",X"19",X"5e",X"23",X"56",X"eb", -- 26e8
  X"c9",X"d1",X"c1",X"c5",X"d5",X"11",X"e0",X"22", -- 26f0
  X"26",X"00",X"69",X"29",X"19",X"5e",X"23",X"56", -- 26f8
  X"eb",X"c9",X"d1",X"c1",X"c5",X"d5",X"11",X"e0", -- 2700
  X"24",X"26",X"00",X"69",X"29",X"19",X"5e",X"23", -- 2708
  X"56",X"eb",X"c9",X"44",X"4d",X"21",X"00",X"00", -- 2710
  X"79",X"0f",X"d2",X"1e",X"27",X"19",X"af",X"78", -- 2718
  X"1f",X"47",X"79",X"1f",X"4f",X"b0",X"c8",X"af", -- 2720
  X"7b",X"17",X"5f",X"7a",X"17",X"57",X"b3",X"c8", -- 2728
  X"c3",X"18",X"27",X"44",X"4d",X"7a",X"a8",X"f5", -- 2730
  X"7a",X"b7",X"fc",X"74",X"27",X"78",X"b7",X"fc", -- 2738
  X"7c",X"27",X"3e",X"10",X"f5",X"eb",X"11",X"00", -- 2740
  X"00",X"29",X"cd",X"84",X"27",X"ca",X"60",X"27", -- 2748
  X"cd",X"8c",X"27",X"fa",X"60",X"27",X"7d",X"f6", -- 2750
  X"01",X"6f",X"7b",X"91",X"5f",X"7a",X"98",X"57", -- 2758
  X"f1",X"3d",X"ca",X"69",X"27",X"f5",X"c3",X"49", -- 2760
  X"27",X"f1",X"f0",X"cd",X"74",X"27",X"eb",X"cd", -- 2768
  X"74",X"27",X"eb",X"c9",X"7a",X"2f",X"57",X"7b", -- 2770
  X"2f",X"5f",X"13",X"c9",X"78",X"2f",X"47",X"79", -- 2778
  X"2f",X"4f",X"03",X"c9",X"7b",X"17",X"5f",X"7a", -- 2780
  X"17",X"57",X"b3",X"c9",X"7b",X"91",X"7a",X"98", -- 2788
  X"c9",X"eb",X"e1",X"4e",X"23",X"46",X"23",X"78", -- 2790
  X"b1",X"ca",X"aa",X"27",X"7e",X"23",X"bb",X"7e", -- 2798
  X"23",X"c2",X"93",X"27",X"ba",X"c2",X"93",X"27", -- 27a0
  X"60",X"69",X"e9",X"eb",X"1d",X"f8",X"7c",X"17", -- 27a8
  X"7c",X"1f",X"67",X"7d",X"1f",X"6f",X"c3",X"ac", -- 27b0
  X"27",X"eb",X"1d",X"f8",X"29",X"c3",X"ba",X"27", -- 27b8
  X"e9",X"19",X"c3",X"c8",X"27",X"23",X"23",X"39", -- 27c0
  X"7e",X"6f",X"07",X"9f",X"67",X"c9",X"19",X"c3", -- 27c8
  X"d5",X"27",X"23",X"23",X"39",X"7e",X"23",X"66", -- 27d0
  X"6f",X"c9",X"23",X"23",X"39",X"54",X"5d",X"cd", -- 27d8
  X"c8",X"27",X"2b",X"7d",X"12",X"c9",X"23",X"23", -- 27e0
  X"39",X"54",X"5d",X"cd",X"c8",X"27",X"23",X"7d", -- 27e8
  X"12",X"c9",X"19",X"c1",X"d1",X"c5",X"7d",X"12", -- 27f0
  X"c9",X"23",X"23",X"39",X"54",X"5d",X"cd",X"d5", -- 27f8
  X"27",X"2b",X"c3",X"15",X"28",X"23",X"23",X"39", -- 2800
  X"54",X"5d",X"cd",X"d5",X"27",X"23",X"c3",X"15", -- 2808
  X"28",X"19",X"c1",X"d1",X"c5",X"7d",X"12",X"13", -- 2810
  X"7c",X"12",X"c9",X"7d",X"b3",X"6f",X"7c",X"b2", -- 2818
  X"67",X"c9",X"7d",X"ab",X"6f",X"7c",X"aa",X"67", -- 2820
  X"c9",X"7d",X"a3",X"6f",X"7c",X"a2",X"67",X"c9", -- 2828
  X"cd",X"56",X"28",X"c8",X"2b",X"c9",X"cd",X"56", -- 2830
  X"28",X"c0",X"2b",X"c9",X"eb",X"cd",X"56",X"28", -- 2838
  X"d8",X"2b",X"c9",X"cd",X"56",X"28",X"c8",X"d8", -- 2840
  X"2b",X"c9",X"cd",X"56",X"28",X"d0",X"2b",X"c9", -- 2848
  X"cd",X"56",X"28",X"d8",X"2b",X"c9",X"7c",X"ee", -- 2850
  X"80",X"67",X"7a",X"ee",X"80",X"bc",X"c2",X"63", -- 2858
  X"28",X"7b",X"bd",X"21",X"01",X"00",X"c9",X"cd", -- 2860
  X"81",X"28",X"d0",X"2b",X"c9",X"cd",X"81",X"28", -- 2868
  X"d8",X"2b",X"c9",X"eb",X"cd",X"81",X"28",X"d8", -- 2870
  X"2b",X"c9",X"cd",X"81",X"28",X"c8",X"d8",X"2b", -- 2878
  X"c9",X"7a",X"bc",X"c2",X"88",X"28",X"7b",X"bd", -- 2880
  X"21",X"01",X"00",X"c9",X"7b",X"95",X"6f",X"7a", -- 2888
  X"9c",X"67",X"c9",X"cd",X"98",X"28",X"23",X"c9", -- 2890
  X"7c",X"2f",X"67",X"7d",X"2f",X"6f",X"c9",X"7c", -- 2898
  X"b5",X"c2",X"a7",X"28",X"2e",X"01",X"c9",X"21", -- 28a0
  X"00",X"00",X"c9",X"00",X"00",X"00",X"00",X"00", -- 28a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2900
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2908
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2910
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2918
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2920
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2928
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2930
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2938
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2940
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2948
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2950
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2958
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2960
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2968
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2970
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2978
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2980
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2988
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2990
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2998
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2aa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2aa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ab0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ab8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ac0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ac8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ad0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ad8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ae0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ae8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2af0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2af8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ba0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ba8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2be0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2be8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ca0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ca8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ce0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ce8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2da0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2da8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2db0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2db8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2de0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2de8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2df0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2df8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ea0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ea8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2eb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2eb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ec0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ec8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ed0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ed8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ee0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ee8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ef0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ef8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fe0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fe8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ff0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ff8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3000
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3008
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3010
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3018
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3020
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3028
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3030
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3038
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3040
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3048
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3050
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3058
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3060
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3068
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3070
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3078
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3080
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3088
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3090
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3098
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3100
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3108
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3110
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3118
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3120
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3128
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3130
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3138
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3140
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3148
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3150
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3158
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3160
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3168
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3170
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3178
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3180
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3188
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3190
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3198
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3200
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3208
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3210
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3218
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3220
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3228
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3230
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3238
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3240
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3248
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3250
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3258
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3260
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3268
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3270
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3278
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3280
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3288
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3290
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3298
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3300
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3308
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3310
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3318
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3320
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3328
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3330
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3338
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3340
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3348
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3350
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3358
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3360
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3368
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3370
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3378
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3380
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3388
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3390
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3398
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3400
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3408
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3410
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3418
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3420
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3428
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3430
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3438
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3440
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3448
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3450
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3458
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3460
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3468
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3470
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3478
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3480
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3488
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3490
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3498
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3500
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3508
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3510
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3518
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3520
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3528
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3530
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3538
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3540
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3548
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3550
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3558
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3560
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3568
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3570
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3578
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3580
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3588
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3590
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3598
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3600
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3608
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3610
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3618
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3620
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3628
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3630
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3638
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3640
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3648
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3650
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3658
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3660
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3668
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3670
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3678
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3680
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3688
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3690
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3698
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3700
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3708
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3710
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3718
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3720
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3728
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3730
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3738
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3740
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3748
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3750
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3758
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3760
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3768
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3770
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3778
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3780
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3788
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3790
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3798
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3800
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3808
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3810
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3818
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3820
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3828
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3830
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3838
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3840
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3848
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3850
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3858
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3860
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3868
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3870
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3878
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3880
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3888
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3890
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3898
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3900
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3908
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3910
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3918
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3920
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3928
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3930
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3938
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3940
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3948
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3950
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3958
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3960
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3968
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3970
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3978
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3980
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3988
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3990
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3998
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3aa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3aa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ab0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ab8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ac0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ac8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ad0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ad8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ae0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ae8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3af0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3af8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ba0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ba8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3be0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3be8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ca0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ca8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ce0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ce8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3da0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3da8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3db0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3db8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3de0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3de8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3df0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3df8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ea0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ea8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3eb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3eb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ec0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ec8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ed0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ed8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ee0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ee8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ef0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ef8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fe0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fe8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ff0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"  -- 3ff8
  );

end package obj_code_pkg;
