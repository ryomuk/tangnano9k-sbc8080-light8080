-------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
-------------------------------------------------------------------------------
-- Generated from "PTBEXSA.BIN"
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Package with utility functions for handling SoC object code.
use work.mcu80_pkg.all;

package obj_code_pkg is

-- Object code initialization constant.
constant object_code : obj_code_t(0 to 16383) := (
  X"c3",X"d4",X"00",X"00",X"00",X"f5",X"79",X"07", -- 0000
  X"81",X"4f",X"f1",X"06",X"00",X"21",X"12",X"00", -- 0008
  X"09",X"e9",X"c3",X"d4",X"00",X"c3",X"7c",X"00", -- 0010
  X"c3",X"ab",X"00",X"c3",X"7c",X"00",X"c3",X"ab", -- 0018
  X"00",X"c3",X"ab",X"00",X"c3",X"c0",X"00",X"db", -- 0020
  X"01",X"e6",X"02",X"ca",X"27",X"00",X"db",X"00", -- 0028
  X"c9",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0030
  X"f3",X"f5",X"c5",X"d5",X"e5",X"cd",X"27",X"00", -- 0038
  X"fe",X"11",X"ca",X"4a",X"00",X"fe",X"13",X"c2", -- 0040
  X"50",X"00",X"32",X"03",X"fe",X"c3",X"76",X"00", -- 0048
  X"57",X"3a",X"00",X"fe",X"fe",X"ff",X"ca",X"76", -- 0050
  X"00",X"fe",X"af",X"c2",X"63",X"00",X"1e",X"13", -- 0058
  X"cd",X"ab",X"00",X"3c",X"32",X"00",X"fe",X"3a", -- 0060
  X"02",X"fe",X"4f",X"06",X"00",X"21",X"04",X"fe", -- 0068
  X"09",X"72",X"3c",X"32",X"02",X"fe",X"e1",X"d1", -- 0070
  X"c1",X"f1",X"fb",X"c9",X"c5",X"d5",X"e5",X"3a", -- 0078
  X"00",X"fe",X"fe",X"00",X"ca",X"7f",X"00",X"f3", -- 0080
  X"fe",X"af",X"c2",X"92",X"00",X"1e",X"11",X"cd", -- 0088
  X"ab",X"00",X"3d",X"32",X"00",X"fe",X"3a",X"01", -- 0090
  X"fe",X"4f",X"06",X"00",X"21",X"04",X"fe",X"09", -- 0098
  X"56",X"3c",X"32",X"01",X"fe",X"7a",X"fb",X"e1", -- 00a0
  X"d1",X"c1",X"c9",X"f5",X"3a",X"03",X"fe",X"fe", -- 00a8
  X"13",X"ca",X"ac",X"00",X"db",X"01",X"e6",X"01", -- 00b0
  X"ca",X"b4",X"00",X"7b",X"d3",X"00",X"f1",X"c9", -- 00b8
  X"f5",X"7b",X"fe",X"ff",X"ca",X"ca",X"00",X"c3", -- 00c0
  X"b4",X"00",X"f1",X"3a",X"00",X"fe",X"fe",X"00", -- 00c8
  X"c8",X"c3",X"7c",X"00",X"31",X"00",X"fe",X"3e", -- 00d0
  X"11",X"32",X"03",X"fe",X"3e",X"00",X"32",X"00", -- 00d8
  X"fe",X"32",X"01",X"fe",X"32",X"02",X"fe",X"d3", -- 00e0
  X"01",X"d3",X"01",X"d3",X"01",X"3e",X"40",X"d3", -- 00e8
  X"01",X"3e",X"4e",X"d3",X"01",X"3e",X"37",X"d3", -- 00f0
  X"01",X"fb",X"c3",X"00",X"01",X"00",X"00",X"00", -- 00f8
  X"31",X"00",X"fe",X"21",X"14",X"90",X"22",X"00", -- 0100
  X"90",X"cd",X"c0",X"08",X"11",X"7e",X"08",X"97", -- 0108
  X"cd",X"b2",X"08",X"11",X"93",X"08",X"97",X"cd", -- 0110
  X"b2",X"08",X"11",X"a2",X"08",X"97",X"cd",X"b2", -- 0118
  X"08",X"cd",X"c0",X"08",X"11",X"6a",X"08",X"97", -- 0120
  X"cd",X"b2",X"08",X"21",X"32",X"01",X"22",X"02", -- 0128
  X"90",X"21",X"00",X"00",X"22",X"08",X"90",X"22", -- 0130
  X"04",X"90",X"3e",X"3e",X"cd",X"9a",X"01",X"d5", -- 0138
  X"11",X"37",X"f0",X"cd",X"ec",X"07",X"cd",X"69", -- 0140
  X"02",X"7c",X"b5",X"c1",X"ca",X"22",X"02",X"1b", -- 0148
  X"7c",X"12",X"1b",X"7d",X"12",X"c5",X"d5",X"79", -- 0150
  X"93",X"f5",X"cd",X"de",X"01",X"d5",X"c2",X"71", -- 0158
  X"01",X"d5",X"cd",X"fc",X"01",X"c1",X"2a",X"00", -- 0160
  X"90",X"cd",X"08",X"02",X"60",X"69",X"22",X"00", -- 0168
  X"90",X"c1",X"2a",X"00",X"90",X"f1",X"e5",X"fe", -- 0170
  X"03",X"ca",X"21",X"01",X"85",X"6f",X"3e",X"00", -- 0178
  X"8c",X"67",X"11",X"00",X"f0",X"cd",X"4d",X"07", -- 0180
  X"d2",X"3b",X"08",X"22",X"00",X"90",X"d1",X"cd", -- 0188
  X"13",X"02",X"d1",X"e1",X"cd",X"08",X"02",X"c3", -- 0190
  X"3a",X"01",X"cd",X"c2",X"08",X"11",X"37",X"f0", -- 0198
  X"cd",X"dd",X"08",X"ca",X"a0",X"01",X"fe",X"0a", -- 01a0
  X"ca",X"a0",X"01",X"b7",X"ca",X"a0",X"01",X"fe", -- 01a8
  X"08",X"ca",X"c7",X"01",X"fe",X"18",X"ca",X"d6", -- 01b0
  X"01",X"cd",X"c2",X"08",X"12",X"13",X"fe",X"0d", -- 01b8
  X"c8",X"7b",X"fe",X"87",X"c2",X"a0",X"01",X"7b", -- 01c0
  X"fe",X"37",X"ca",X"a0",X"01",X"1b",X"3e",X"08", -- 01c8
  X"cd",X"c2",X"08",X"c3",X"a0",X"01",X"cd",X"c0", -- 01d0
  X"08",X"3e",X"40",X"c3",X"9a",X"01",X"7c",X"b7", -- 01d8
  X"fa",X"34",X"08",X"11",X"14",X"90",X"e5",X"2a", -- 01e0
  X"00",X"90",X"2b",X"cd",X"4d",X"07",X"e1",X"d8", -- 01e8
  X"1a",X"95",X"47",X"13",X"1a",X"9c",X"da",X"fd", -- 01f0
  X"01",X"1b",X"b0",X"c9",X"13",X"13",X"1a",X"fe", -- 01f8
  X"0d",X"c2",X"fd",X"01",X"13",X"c3",X"e6",X"01", -- 0200
  X"cd",X"4d",X"07",X"c8",X"1a",X"02",X"13",X"03", -- 0208
  X"c3",X"08",X"02",X"78",X"92",X"c2",X"1b",X"02", -- 0210
  X"79",X"93",X"c8",X"1b",X"2b",X"1a",X"77",X"c3", -- 0218
  X"13",X"02",X"21",X"70",X"02",X"cd",X"69",X"02", -- 0220
  X"d5",X"1a",X"13",X"fe",X"2e",X"ca",X"46",X"02", -- 0228
  X"23",X"be",X"ca",X"29",X"02",X"3e",X"7f",X"1b", -- 0230
  X"be",X"da",X"4d",X"02",X"23",X"be",X"d2",X"3c", -- 0238
  X"02",X"23",X"d1",X"c3",X"28",X"02",X"3e",X"7f", -- 0240
  X"23",X"be",X"d2",X"48",X"02",X"7e",X"23",X"6e", -- 0248
  X"e6",X"7f",X"67",X"f1",X"e9",X"e3",X"cd",X"69", -- 0250
  X"02",X"be",X"23",X"ca",X"65",X"02",X"c5",X"4e", -- 0258
  X"06",X"00",X"09",X"c1",X"1b",X"13",X"23",X"e3", -- 0260
  X"c9",X"1a",X"fe",X"20",X"c0",X"13",X"c3",X"69", -- 0268
  X"02",X"4c",X"49",X"53",X"54",X"84",X"62",X"52", -- 0270
  X"55",X"4e",X"85",X"df",X"4e",X"45",X"57",X"82", -- 0278
  X"f0",X"53",X"59",X"53",X"54",X"45",X"4d",X"82", -- 0280
  X"ff",X"4d",X"4f",X"4e",X"82",X"d8",X"4e",X"45", -- 0288
  X"58",X"54",X"83",X"b4",X"4c",X"45",X"54",X"85", -- 0290
  X"ad",X"49",X"4e",X"50",X"55",X"54",X"85",X"51", -- 0298
  X"49",X"46",X"84",X"4e",X"47",X"4f",X"54",X"4f", -- 02a0
  X"85",X"ce",X"47",X"4f",X"53",X"55",X"42",X"83", -- 02a8
  X"04",X"52",X"45",X"54",X"55",X"52",X"4e",X"83", -- 02b0
  X"26",X"52",X"45",X"4d",X"84",X"56",X"46",X"4f", -- 02b8
  X"52",X"83",X"41",X"50",X"52",X"49",X"4e",X"54", -- 02c0
  X"84",X"8f",X"53",X"54",X"4f",X"50",X"82",X"f9", -- 02c8
  X"45",X"58",X"45",X"43",X"82",X"db",X"85",X"a5", -- 02d0
  X"c3",X"00",X"09",X"cd",X"20",X"06",X"f5",X"c5", -- 02d8
  X"d5",X"11",X"ea",X"02",X"d5",X"11",X"00",X"80", -- 02e0
  X"19",X"e9",X"d1",X"c1",X"f1",X"c3",X"fe",X"05", -- 02e8
  X"cd",X"17",X"06",X"21",X"14",X"90",X"22",X"00", -- 02f0
  X"90",X"cd",X"17",X"06",X"c3",X"21",X"01",X"0e", -- 02f8
  X"00",X"cd",X"05",X"00",X"cd",X"09",X"04",X"cd", -- 0300
  X"20",X"06",X"d5",X"cd",X"de",X"01",X"c2",X"35", -- 0308
  X"08",X"2a",X"02",X"90",X"e5",X"2a",X"04",X"90", -- 0310
  X"e5",X"21",X"00",X"00",X"22",X"08",X"90",X"39", -- 0318
  X"22",X"04",X"90",X"c3",X"ee",X"05",X"cd",X"17", -- 0320
  X"06",X"2a",X"04",X"90",X"7c",X"b5",X"ca",X"2d", -- 0328
  X"08",X"f9",X"e1",X"22",X"04",X"90",X"e1",X"22", -- 0330
  X"02",X"90",X"d1",X"cd",X"32",X"04",X"c3",X"fe", -- 0338
  X"05",X"cd",X"09",X"04",X"cd",X"b8",X"05",X"2b", -- 0340
  X"22",X"08",X"90",X"21",X"50",X"03",X"c3",X"25", -- 0348
  X"02",X"54",X"4f",X"83",X"57",X"88",X"2d",X"cd", -- 0350
  X"20",X"06",X"22",X"0c",X"90",X"21",X"62",X"03", -- 0358
  X"c3",X"25",X"02",X"53",X"54",X"45",X"50",X"83", -- 0360
  X"6b",X"83",X"71",X"cd",X"20",X"06",X"c3",X"74", -- 0368
  X"03",X"21",X"01",X"00",X"22",X"0a",X"90",X"2a", -- 0370
  X"02",X"90",X"22",X"0e",X"90",X"eb",X"22",X"10", -- 0378
  X"90",X"01",X"0a",X"00",X"2a",X"08",X"90",X"eb", -- 0380
  X"60",X"68",X"39",X"3e",X"09",X"7e",X"23",X"b6", -- 0388
  X"ca",X"ad",X"03",X"7e",X"2b",X"ba",X"c2",X"8c", -- 0390
  X"03",X"7e",X"bb",X"c2",X"8c",X"03",X"eb",X"21", -- 0398
  X"00",X"00",X"39",X"44",X"4d",X"21",X"0a",X"00", -- 03a0
  X"19",X"cd",X"13",X"02",X"f9",X"2a",X"10",X"90", -- 03a8
  X"eb",X"c3",X"fe",X"05",X"cd",X"b8",X"07",X"da", -- 03b0
  X"2d",X"08",X"22",X"06",X"90",X"d5",X"eb",X"2a", -- 03b8
  X"08",X"90",X"7c",X"b5",X"ca",X"2e",X"08",X"cd", -- 03c0
  X"4d",X"07",X"ca",X"d7",X"03",X"d1",X"cd",X"32", -- 03c8
  X"04",X"2a",X"06",X"90",X"c3",X"bd",X"03",X"5e", -- 03d0
  X"23",X"56",X"2a",X"0a",X"90",X"e5",X"19",X"eb", -- 03d8
  X"2a",X"08",X"90",X"73",X"23",X"72",X"2a",X"0c", -- 03e0
  X"90",X"f1",X"b7",X"f2",X"ef",X"03",X"eb",X"cd", -- 03e8
  X"47",X"07",X"d1",X"da",X"03",X"04",X"2a",X"0e", -- 03f0
  X"90",X"22",X"02",X"90",X"2a",X"10",X"90",X"eb", -- 03f8
  X"c3",X"fe",X"05",X"cd",X"32",X"04",X"c3",X"fe", -- 0400
  X"05",X"21",X"a5",X"f0",X"cd",X"3b",X"07",X"c1", -- 0408
  X"39",X"d2",X"3b",X"08",X"2a",X"08",X"90",X"7c", -- 0410
  X"b5",X"ca",X"2f",X"04",X"2a",X"10",X"90",X"e5", -- 0418
  X"2a",X"0e",X"90",X"e5",X"2a",X"0c",X"90",X"e5", -- 0420
  X"2a",X"0a",X"90",X"e5",X"2a",X"08",X"90",X"e5", -- 0428
  X"c5",X"c9",X"c1",X"e1",X"22",X"08",X"90",X"7c", -- 0430
  X"b5",X"ca",X"4c",X"04",X"e1",X"22",X"0a",X"90", -- 0438
  X"e1",X"22",X"0c",X"90",X"e1",X"22",X"0e",X"90", -- 0440
  X"e1",X"22",X"10",X"90",X"c5",X"c9",X"cd",X"20", -- 0448
  X"06",X"7c",X"b5",X"c2",X"f5",X"05",X"21",X"00", -- 0450
  X"00",X"cd",X"fe",X"01",X"d2",X"ee",X"05",X"c3", -- 0458
  X"21",X"01",X"cd",X"ec",X"07",X"cd",X"17",X"06", -- 0460
  X"cd",X"de",X"01",X"da",X"21",X"01",X"cd",X"7a", -- 0468
  X"04",X"cd",X"dd",X"08",X"cd",X"e6",X"01",X"c3", -- 0470
  X"6b",X"04",X"1a",X"6f",X"13",X"1a",X"67",X"13", -- 0478
  X"0e",X"04",X"cd",X"05",X"05",X"3e",X"20",X"cd", -- 0480
  X"c2",X"08",X"97",X"cd",X"b2",X"08",X"c9",X"0e", -- 0488
  X"06",X"cd",X"55",X"02",X"3b",X"06",X"cd",X"c0", -- 0490
  X"08",X"c3",X"f5",X"05",X"cd",X"55",X"02",X"0d", -- 0498
  X"06",X"cd",X"c0",X"08",X"c3",X"e5",X"05",X"cd", -- 04a0
  X"55",X"02",X"23",X"07",X"cd",X"20",X"06",X"4d", -- 04a8
  X"c3",X"b9",X"04",X"cd",X"d5",X"04",X"c3",X"ca", -- 04b0
  X"04",X"cd",X"55",X"02",X"2c",X"06",X"cd",X"04", -- 04b8
  X"06",X"c3",X"a7",X"04",X"cd",X"c0",X"08",X"c3", -- 04c0
  X"fe",X"05",X"cd",X"20",X"06",X"c5",X"cd",X"05", -- 04c8
  X"05",X"c1",X"c3",X"b9",X"04",X"cd",X"55",X"02", -- 04d0
  X"22",X"05",X"3e",X"22",X"c3",X"e6",X"04",X"cd", -- 04d8
  X"55",X"02",X"27",X"0e",X"3e",X"27",X"cd",X"b2", -- 04e0
  X"08",X"fe",X"0d",X"e1",X"ca",X"e5",X"05",X"c3", -- 04e8
  X"00",X"05",X"cd",X"55",X"02",X"5f",X"0d",X"3e", -- 04f0
  X"8d",X"cd",X"c2",X"08",X"cd",X"c2",X"08",X"e1", -- 04f8
  X"23",X"23",X"23",X"e9",X"c9",X"d5",X"11",X"0a", -- 0500
  X"00",X"d5",X"42",X"0d",X"cd",X"38",X"07",X"f2", -- 0508
  X"15",X"05",X"06",X"2d",X"0d",X"c5",X"cd",X"1b", -- 0510
  X"07",X"78",X"b1",X"ca",X"26",X"05",X"e3",X"2d", -- 0518
  X"e5",X"60",X"69",X"c3",X"16",X"05",X"c1",X"0d", -- 0520
  X"79",X"b7",X"fa",X"35",X"05",X"3e",X"20",X"cd", -- 0528
  X"c2",X"08",X"c3",X"27",X"05",X"78",X"cd",X"c2", -- 0530
  X"08",X"5d",X"7b",X"fe",X"0a",X"d1",X"c8",X"c6", -- 0538
  X"30",X"cd",X"c2",X"08",X"c3",X"3a",X"05",X"2a", -- 0540
  X"06",X"90",X"f9",X"e1",X"22",X"02",X"90",X"d1", -- 0548
  X"d1",X"d5",X"cd",X"d5",X"04",X"c3",X"61",X"05", -- 0550
  X"cd",X"b8",X"07",X"da",X"9c",X"05",X"c3",X"73", -- 0558
  X"05",X"d5",X"cd",X"b8",X"07",X"da",X"2d",X"08", -- 0560
  X"1a",X"4f",X"97",X"12",X"d1",X"cd",X"b2",X"08", -- 0568
  X"79",X"1b",X"12",X"d5",X"eb",X"2a",X"02",X"90", -- 0570
  X"e5",X"21",X"51",X"05",X"22",X"02",X"90",X"21", -- 0578
  X"00",X"00",X"39",X"22",X"06",X"90",X"d5",X"3e", -- 0580
  X"3a",X"cd",X"9a",X"01",X"11",X"37",X"f0",X"cd", -- 0588
  X"20",X"06",X"d1",X"eb",X"73",X"23",X"72",X"e1", -- 0590
  X"22",X"02",X"90",X"d1",X"f1",X"cd",X"55",X"02", -- 0598
  X"2c",X"5c",X"c3",X"51",X"05",X"cd",X"0d",X"06", -- 05a0
  X"fe",X"0d",X"ca",X"fe",X"05",X"cd",X"b8",X"05", -- 05a8
  X"cd",X"55",X"02",X"2c",X"49",X"c3",X"ad",X"05", -- 05b0
  X"cd",X"b8",X"07",X"da",X"2d",X"08",X"e5",X"cd", -- 05b8
  X"55",X"02",X"3d",X"3d",X"cd",X"20",X"06",X"44", -- 05c0
  X"4d",X"e1",X"71",X"23",X"70",X"c9",X"cd",X"20", -- 05c8
  X"06",X"d5",X"cd",X"17",X"06",X"cd",X"de",X"01", -- 05d0
  X"c2",X"35",X"08",X"f1",X"c3",X"ee",X"05",X"cd", -- 05d8
  X"17",X"06",X"11",X"14",X"90",X"21",X"00",X"00", -- 05e0
  X"cd",X"e6",X"01",X"da",X"21",X"01",X"eb",X"22", -- 05e8
  X"02",X"90",X"eb",X"13",X"13",X"cd",X"dd",X"08", -- 05f0
  X"21",X"8d",X"02",X"c3",X"25",X"02",X"cd",X"04", -- 05f8
  X"06",X"c3",X"2d",X"08",X"cd",X"55",X"02",X"3b", -- 0600
  X"04",X"f1",X"c3",X"f5",X"05",X"cd",X"55",X"02", -- 0608
  X"0d",X"04",X"f1",X"c3",X"e5",X"05",X"c9",X"cd", -- 0610
  X"69",X"02",X"fe",X"0d",X"c8",X"c3",X"2d",X"08", -- 0618
  X"cd",X"7f",X"06",X"e5",X"21",X"29",X"06",X"c3", -- 0620
  X"25",X"02",X"3e",X"3d",X"86",X"41",X"3c",X"3e", -- 0628
  X"86",X"47",X"3e",X"86",X"4d",X"3d",X"86",X"5c", -- 0630
  X"3c",X"3d",X"86",X"54",X"3c",X"86",X"62",X"86", -- 0638
  X"68",X"cd",X"6a",X"06",X"d8",X"6f",X"c9",X"cd", -- 0640
  X"6a",X"06",X"c8",X"6f",X"c9",X"cd",X"6a",X"06", -- 0648
  X"c8",X"d8",X"6f",X"c9",X"cd",X"6a",X"06",X"6f", -- 0650
  X"c8",X"d8",X"6c",X"c9",X"cd",X"6a",X"06",X"c0", -- 0658
  X"6f",X"c9",X"cd",X"6a",X"06",X"d0",X"6f",X"c9", -- 0660
  X"e1",X"c9",X"79",X"e1",X"c1",X"e5",X"c5",X"4f", -- 0668
  X"cd",X"7f",X"06",X"eb",X"e3",X"cd",X"47",X"07", -- 0670
  X"d1",X"21",X"00",X"00",X"3e",X"01",X"c9",X"cd", -- 0678
  X"55",X"02",X"2d",X"06",X"21",X"00",X"00",X"c3", -- 0680
  X"a3",X"06",X"cd",X"55",X"02",X"2b",X"00",X"cd", -- 0688
  X"bb",X"06",X"cd",X"55",X"02",X"2b",X"07",X"e5", -- 0690
  X"cd",X"bb",X"06",X"c3",X"aa",X"06",X"cd",X"55", -- 0698
  X"02",X"2d",X"8d",X"e5",X"cd",X"bb",X"06",X"cd", -- 06a0
  X"3b",X"07",X"eb",X"e3",X"7c",X"aa",X"7a",X"19", -- 06a8
  X"d1",X"fa",X"92",X"06",X"ac",X"f2",X"92",X"06", -- 06b0
  X"c3",X"34",X"08",X"cd",X"53",X"07",X"cd",X"55", -- 06b8
  X"02",X"2a",X"2b",X"e5",X"cd",X"53",X"07",X"06", -- 06c0
  X"00",X"cd",X"38",X"07",X"eb",X"e3",X"cd",X"38", -- 06c8
  X"07",X"7c",X"b7",X"ca",X"dc",X"06",X"7a",X"b2", -- 06d0
  X"eb",X"c2",X"35",X"08",X"7d",X"2e",X"00",X"b7", -- 06d8
  X"ca",X"0d",X"07",X"19",X"da",X"35",X"08",X"3d", -- 06e0
  X"c2",X"e3",X"06",X"c3",X"0d",X"07",X"cd",X"55", -- 06e8
  X"02",X"2f",X"3d",X"e5",X"cd",X"53",X"07",X"06", -- 06f0
  X"00",X"cd",X"38",X"07",X"eb",X"e3",X"cd",X"38", -- 06f8
  X"07",X"7a",X"b3",X"ca",X"35",X"08",X"c5",X"cd", -- 0700
  X"1b",X"07",X"60",X"69",X"c1",X"d1",X"7c",X"b7", -- 0708
  X"fa",X"34",X"08",X"78",X"b7",X"fc",X"3b",X"07", -- 0710
  X"c3",X"be",X"06",X"e5",X"6c",X"26",X"00",X"cd", -- 0718
  X"26",X"07",X"41",X"7d",X"e1",X"67",X"0e",X"ff", -- 0720
  X"0c",X"cd",X"31",X"07",X"d2",X"28",X"07",X"19", -- 0728
  X"c9",X"7d",X"93",X"6f",X"7c",X"9a",X"67",X"c9", -- 0730
  X"7c",X"b7",X"f0",X"7c",X"2f",X"67",X"7d",X"2f", -- 0738
  X"6f",X"23",X"78",X"ee",X"80",X"47",X"c9",X"7c", -- 0740
  X"aa",X"f2",X"4d",X"07",X"eb",X"7c",X"ba",X"c0", -- 0748
  X"7d",X"bb",X"c9",X"21",X"58",X"07",X"c3",X"25", -- 0750
  X"02",X"52",X"4e",X"44",X"87",X"6b",X"41",X"42", -- 0758
  X"53",X"87",X"94",X"53",X"49",X"5a",X"45",X"87", -- 0760
  X"a0",X"87",X"ad",X"cd",X"1f",X"08",X"7c",X"b7", -- 0768
  X"fa",X"34",X"08",X"b5",X"ca",X"34",X"08",X"d5", -- 0770
  X"e5",X"2a",X"12",X"90",X"7c",X"e6",X"07",X"67", -- 0778
  X"11",X"00",X"01",X"19",X"5e",X"23",X"56",X"22", -- 0780
  X"12",X"90",X"e1",X"eb",X"c5",X"cd",X"1b",X"07", -- 0788
  X"c1",X"d1",X"23",X"c9",X"cd",X"1f",X"08",X"cd", -- 0790
  X"38",X"07",X"7c",X"b4",X"fa",X"34",X"08",X"c9", -- 0798
  X"2a",X"00",X"90",X"d5",X"eb",X"21",X"00",X"f0", -- 07a0
  X"cd",X"31",X"07",X"d1",X"c9",X"cd",X"b8",X"07", -- 07a8
  X"da",X"19",X"08",X"7e",X"23",X"66",X"6f",X"c9", -- 07b0
  X"cd",X"69",X"02",X"d6",X"40",X"d8",X"c2",X"dc", -- 07b8
  X"07",X"13",X"cd",X"1f",X"08",X"29",X"da",X"34", -- 07c0
  X"08",X"d5",X"eb",X"cd",X"a0",X"07",X"cd",X"4d", -- 07c8
  X"07",X"da",X"3c",X"08",X"21",X"00",X"f0",X"cd", -- 07d0
  X"31",X"07",X"d1",X"c9",X"fe",X"1b",X"3f",X"d8", -- 07d8
  X"13",X"21",X"00",X"f0",X"07",X"85",X"6f",X"3e", -- 07e0
  X"00",X"8c",X"67",X"c9",X"21",X"00",X"00",X"44", -- 07e8
  X"cd",X"69",X"02",X"fe",X"30",X"d8",X"fe",X"3a", -- 07f0
  X"d0",X"3e",X"f0",X"a4",X"c2",X"34",X"08",X"04", -- 07f8
  X"c5",X"44",X"4d",X"29",X"29",X"09",X"29",X"1a", -- 0800
  X"13",X"e6",X"0f",X"85",X"6f",X"3e",X"00",X"8c", -- 0808
  X"67",X"c1",X"1a",X"fa",X"34",X"08",X"c3",X"f3", -- 0810
  X"07",X"cd",X"ec",X"07",X"78",X"b7",X"c0",X"cd", -- 0818
  X"55",X"02",X"28",X"09",X"cd",X"20",X"06",X"cd", -- 0820
  X"55",X"02",X"29",X"01",X"c9",X"d5",X"11",X"72", -- 0828
  X"08",X"c3",X"3f",X"08",X"d5",X"11",X"6d",X"08", -- 0830
  X"c3",X"3f",X"08",X"d5",X"11",X"78",X"08",X"97", -- 0838
  X"cd",X"b2",X"08",X"d1",X"1a",X"f5",X"97",X"12", -- 0840
  X"2a",X"02",X"90",X"e5",X"7e",X"23",X"b6",X"d1", -- 0848
  X"ca",X"21",X"01",X"7e",X"b7",X"fa",X"47",X"05", -- 0850
  X"cd",X"7a",X"04",X"1b",X"f1",X"12",X"3e",X"3f", -- 0858
  X"cd",X"c2",X"08",X"97",X"cd",X"b2",X"08",X"c3", -- 0860
  X"21",X"01",X"4f",X"4b",X"0d",X"48",X"4f",X"57", -- 0868
  X"3f",X"0d",X"57",X"48",X"41",X"54",X"3f",X"0d", -- 0870
  X"53",X"4f",X"52",X"52",X"59",X"0d",X"50",X"41", -- 0878
  X"4c",X"4f",X"20",X"41",X"4c",X"54",X"4f",X"20", -- 0880
  X"54",X"49",X"4e",X"59",X"20",X"42",X"41",X"53", -- 0888
  X"49",X"43",X"0d",X"4d",X"4f",X"4e",X"38",X"30", -- 0890
  X"20",X"45",X"58",X"54",X"45",X"4e",X"44",X"45", -- 0898
  X"44",X"0d",X"53",X"42",X"43",X"38",X"30",X"38", -- 08a0
  X"30",X"20",X"45",X"44",X"49",X"54",X"49",X"4f", -- 08a8
  X"4e",X"0d",X"47",X"1a",X"13",X"b8",X"c8",X"cd", -- 08b0
  X"c2",X"08",X"fe",X"0d",X"c2",X"b3",X"08",X"c9", -- 08b8
  X"3e",X"0d",X"f5",X"c5",X"d5",X"e5",X"0e",X"02", -- 08c0
  X"e6",X"7f",X"5f",X"cd",X"05",X"00",X"e1",X"d1", -- 08c8
  X"c1",X"f1",X"fe",X"0d",X"c0",X"3e",X"0a",X"cd", -- 08d0
  X"c2",X"08",X"3e",X"0d",X"c9",X"c5",X"d5",X"e5", -- 08d8
  X"0e",X"06",X"1e",X"ff",X"cd",X"05",X"00",X"e1", -- 08e0
  X"d1",X"c1",X"e6",X"7f",X"c8",X"fe",X"1b",X"c2", -- 08e8
  X"f7",X"08",X"33",X"33",X"c3",X"21",X"01",X"fe", -- 08f0
  X"61",X"d8",X"fe",X"7b",X"d0",X"e6",X"df",X"c9", -- 08f8
  X"21",X"1c",X"fe",X"39",X"f9",X"21",X"e2",X"01", -- 0900
  X"39",X"eb",X"21",X"00",X"80",X"cd",X"8d",X"2f", -- 0908
  X"21",X"90",X"01",X"39",X"e5",X"21",X"42",X"01", -- 0910
  X"39",X"e5",X"21",X"f4",X"00",X"39",X"e5",X"21", -- 0918
  X"a6",X"00",X"39",X"e5",X"21",X"58",X"00",X"39", -- 0920
  X"e5",X"21",X"0a",X"00",X"39",X"eb",X"21",X"00", -- 0928
  X"00",X"7d",X"12",X"d1",X"7d",X"12",X"d1",X"7d", -- 0930
  X"12",X"d1",X"7d",X"12",X"d1",X"7d",X"12",X"d1", -- 0938
  X"7d",X"12",X"21",X"e2",X"01",X"39",X"cd",X"4d", -- 0940
  X"2f",X"e5",X"3e",X"01",X"cd",X"0f",X"19",X"c1", -- 0948
  X"21",X"90",X"01",X"39",X"e5",X"21",X"49",X"00", -- 0950
  X"e5",X"3e",X"02",X"cd",X"90",X"25",X"c1",X"c1", -- 0958
  X"21",X"90",X"01",X"39",X"e5",X"21",X"42",X"01", -- 0960
  X"39",X"e5",X"21",X"a4",X"00",X"39",X"e5",X"3e", -- 0968
  X"03",X"cd",X"2f",X"19",X"c1",X"c1",X"c1",X"21", -- 0970
  X"a0",X"00",X"39",X"e5",X"21",X"52",X"00",X"39", -- 0978
  X"e5",X"21",X"04",X"00",X"39",X"e5",X"3e",X"03", -- 0980
  X"cd",X"ae",X"1a",X"c1",X"c1",X"c1",X"21",X"90", -- 0988
  X"01",X"39",X"cd",X"40",X"2f",X"7c",X"b5",X"ca", -- 0990
  X"ab",X"09",X"21",X"f0",X"00",X"39",X"e5",X"21", -- 0998
  X"42",X"01",X"39",X"e5",X"3e",X"02",X"cd",X"a1", -- 09a0
  X"1e",X"c1",X"c1",X"21",X"f0",X"00",X"39",X"e5", -- 09a8
  X"21",X"09",X"0c",X"e5",X"3e",X"02",X"cd",X"cd", -- 09b0
  X"1e",X"c1",X"c1",X"7c",X"b5",X"c2",X"42",X"0a", -- 09b8
  X"21",X"50",X"00",X"39",X"e5",X"3e",X"01",X"cd", -- 09c0
  X"80",X"1d",X"c1",X"7c",X"b5",X"ca",X"e4",X"09", -- 09c8
  X"21",X"e2",X"01",X"39",X"e5",X"21",X"52",X"00", -- 09d0
  X"39",X"e5",X"3e",X"01",X"cd",X"9b",X"22",X"c1", -- 09d8
  X"d1",X"cd",X"8d",X"2f",X"21",X"00",X"00",X"39", -- 09e0
  X"e5",X"3e",X"01",X"cd",X"80",X"1d",X"c1",X"7c", -- 09e8
  X"b5",X"ca",X"0b",X"0a",X"21",X"e0",X"01",X"39", -- 09f0
  X"e5",X"21",X"02",X"00",X"39",X"e5",X"3e",X"01", -- 09f8
  X"cd",X"9b",X"22",X"c1",X"d1",X"cd",X"8d",X"2f", -- 0a00
  X"c3",X"1f",X"0a",X"21",X"e0",X"01",X"39",X"e5", -- 0a08
  X"21",X"e4",X"01",X"39",X"cd",X"4d",X"2f",X"11", -- 0a10
  X"10",X"00",X"19",X"d1",X"cd",X"8d",X"2f",X"21", -- 0a18
  X"e2",X"01",X"39",X"e5",X"21",X"e4",X"01",X"39", -- 0a20
  X"cd",X"4d",X"2f",X"e5",X"21",X"e4",X"01",X"39", -- 0a28
  X"cd",X"4d",X"2f",X"e5",X"3e",X"02",X"cd",X"32", -- 0a30
  X"0c",X"c1",X"c1",X"d1",X"cd",X"8d",X"2f",X"c3", -- 0a38
  X"00",X"0c",X"21",X"f0",X"00",X"39",X"e5",X"21", -- 0a40
  X"0e",X"0c",X"e5",X"3e",X"02",X"cd",X"cd",X"1e", -- 0a48
  X"c1",X"c1",X"7c",X"b5",X"c2",X"d4",X"0a",X"21", -- 0a50
  X"50",X"00",X"39",X"e5",X"3e",X"01",X"cd",X"80", -- 0a58
  X"1d",X"c1",X"7c",X"b5",X"ca",X"7b",X"0a",X"21", -- 0a60
  X"e2",X"01",X"39",X"e5",X"21",X"52",X"00",X"39", -- 0a68
  X"e5",X"3e",X"01",X"cd",X"9b",X"22",X"c1",X"d1", -- 0a70
  X"cd",X"8d",X"2f",X"21",X"00",X"00",X"39",X"e5", -- 0a78
  X"3e",X"01",X"cd",X"80",X"1d",X"c1",X"7c",X"b5", -- 0a80
  X"ca",X"a2",X"0a",X"21",X"e0",X"01",X"39",X"e5", -- 0a88
  X"21",X"02",X"00",X"39",X"e5",X"3e",X"01",X"cd", -- 0a90
  X"9b",X"22",X"c1",X"d1",X"cd",X"8d",X"2f",X"c3", -- 0a98
  X"b1",X"0a",X"21",X"e0",X"01",X"39",X"eb",X"21", -- 0aa0
  X"e2",X"01",X"39",X"cd",X"4d",X"2f",X"cd",X"8d", -- 0aa8
  X"2f",X"21",X"e2",X"01",X"39",X"e5",X"21",X"e4", -- 0ab0
  X"01",X"39",X"cd",X"4d",X"2f",X"e5",X"21",X"e4", -- 0ab8
  X"01",X"39",X"cd",X"4d",X"2f",X"e5",X"3e",X"02", -- 0ac0
  X"cd",X"83",X"0e",X"c1",X"c1",X"d1",X"cd",X"8d", -- 0ac8
  X"2f",X"c3",X"00",X"0c",X"21",X"40",X"01",X"39", -- 0ad0
  X"cd",X"40",X"2f",X"7c",X"b5",X"c2",X"e3",X"0a", -- 0ad8
  X"c3",X"00",X"0c",X"21",X"40",X"01",X"39",X"e5", -- 0ae0
  X"21",X"13",X"0c",X"e5",X"3e",X"02",X"cd",X"cd", -- 0ae8
  X"1e",X"c1",X"c1",X"7c",X"b5",X"c2",X"ff",X"0a", -- 0af0
  X"af",X"cd",X"dd",X"26",X"c3",X"00",X"0c",X"21", -- 0af8
  X"40",X"01",X"39",X"e5",X"21",X"1a",X"0c",X"e5", -- 0b00
  X"3e",X"02",X"cd",X"cd",X"1e",X"c1",X"c1",X"7c", -- 0b08
  X"b5",X"c2",X"22",X"0b",X"21",X"a0",X"00",X"39", -- 0b10
  X"e5",X"3e",X"01",X"cd",X"7e",X"11",X"c1",X"c3", -- 0b18
  X"00",X"0c",X"21",X"40",X"01",X"39",X"e5",X"21", -- 0b20
  X"1f",X"0c",X"e5",X"3e",X"02",X"cd",X"cd",X"1e", -- 0b28
  X"c1",X"c1",X"7c",X"b5",X"c2",X"78",X"0b",X"21", -- 0b30
  X"50",X"00",X"39",X"e5",X"3e",X"01",X"cd",X"80", -- 0b38
  X"1d",X"c1",X"7c",X"b5",X"ca",X"5c",X"0b",X"21", -- 0b40
  X"50",X"00",X"39",X"e5",X"3e",X"01",X"cd",X"9b", -- 0b48
  X"22",X"c1",X"e5",X"3e",X"01",X"cd",X"ac",X"26", -- 0b50
  X"c1",X"c3",X"75",X"0b",X"21",X"24",X"0c",X"e5", -- 0b58
  X"3e",X"01",X"cd",X"68",X"25",X"c1",X"21",X"50", -- 0b60
  X"00",X"39",X"e5",X"3e",X"01",X"cd",X"68",X"25", -- 0b68
  X"c1",X"af",X"cd",X"d5",X"23",X"c3",X"00",X"0c", -- 0b70
  X"21",X"40",X"01",X"39",X"e5",X"21",X"2b",X"0c", -- 0b78
  X"e5",X"3e",X"02",X"cd",X"cd",X"1e",X"c1",X"c1", -- 0b80
  X"7c",X"b5",X"c2",X"ad",X"0b",X"21",X"e2",X"01", -- 0b88
  X"39",X"e5",X"21",X"e4",X"01",X"39",X"cd",X"4d", -- 0b90
  X"2f",X"e5",X"21",X"a4",X"00",X"39",X"e5",X"3e", -- 0b98
  X"02",X"cd",X"6d",X"10",X"c1",X"c1",X"d1",X"cd", -- 0ba0
  X"8d",X"2f",X"c3",X"00",X"0c",X"21",X"40",X"01", -- 0ba8
  X"39",X"e5",X"3e",X"01",X"cd",X"80",X"1d",X"c1", -- 0bb0
  X"7c",X"b5",X"ca",X"d4",X"0b",X"21",X"e2",X"01", -- 0bb8
  X"39",X"e5",X"21",X"42",X"01",X"39",X"e5",X"3e", -- 0bc0
  X"01",X"cd",X"9b",X"22",X"c1",X"d1",X"cd",X"8d", -- 0bc8
  X"2f",X"c3",X"00",X"0c",X"21",X"e2",X"01",X"39", -- 0bd0
  X"e5",X"21",X"e4",X"01",X"39",X"cd",X"4d",X"2f", -- 0bd8
  X"e5",X"21",X"44",X"01",X"39",X"e5",X"21",X"56", -- 0be0
  X"00",X"39",X"e5",X"21",X"08",X"00",X"39",X"e5", -- 0be8
  X"3e",X"04",X"cd",X"ce",X"15",X"eb",X"21",X"08", -- 0bf0
  X"00",X"39",X"f9",X"eb",X"d1",X"cd",X"8d",X"2f", -- 0bf8
  X"c3",X"42",X"09",X"21",X"e4",X"01",X"39",X"f9", -- 0c00
  X"c9",X"4c",X"49",X"53",X"54",X"00",X"44",X"55", -- 0c08
  X"4d",X"50",X"00",X"53",X"59",X"53",X"54",X"45", -- 0c10
  X"4d",X"00",X"48",X"45",X"4c",X"50",X"00",X"45", -- 0c18
  X"58",X"45",X"43",X"00",X"45",X"52",X"52",X"4f", -- 0c20
  X"52",X"2d",X"00",X"44",X"45",X"46",X"49",X"4e", -- 0c28
  X"45",X"00",X"21",X"04",X"00",X"39",X"e5",X"21", -- 0c30
  X"06",X"00",X"39",X"cd",X"4d",X"2f",X"e5",X"3e", -- 0c38
  X"01",X"cd",X"68",X"0c",X"c1",X"d1",X"cd",X"8d", -- 0c40
  X"2f",X"21",X"04",X"00",X"39",X"cd",X"4d",X"2f", -- 0c48
  X"eb",X"c1",X"e1",X"e5",X"c5",X"cd",X"f2",X"2f", -- 0c50
  X"7c",X"b5",X"ca",X"60",X"0c",X"c3",X"32",X"0c", -- 0c58
  X"21",X"04",X"00",X"39",X"cd",X"4d",X"2f",X"c9", -- 0c60
  X"3b",X"c5",X"21",X"20",X"00",X"e5",X"3e",X"01", -- 0c68
  X"cd",X"b7",X"26",X"c1",X"21",X"05",X"00",X"39", -- 0c70
  X"cd",X"4d",X"2f",X"e5",X"3e",X"01",X"cd",X"e3", -- 0c78
  X"23",X"c1",X"21",X"20",X"00",X"e5",X"3e",X"01", -- 0c80
  X"cd",X"b7",X"26",X"c1",X"21",X"02",X"00",X"39", -- 0c88
  X"e5",X"21",X"07",X"00",X"39",X"54",X"5d",X"cd", -- 0c90
  X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"cd", -- 0c98
  X"40",X"2f",X"d1",X"7d",X"12",X"21",X"02",X"00", -- 0ca0
  X"39",X"cd",X"40",X"2f",X"e5",X"3e",X"01",X"cd", -- 0ca8
  X"58",X"2e",X"c1",X"e5",X"3e",X"01",X"cd",X"68", -- 0cb0
  X"25",X"c1",X"21",X"00",X"00",X"39",X"eb",X"21", -- 0cb8
  X"05",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"8d", -- 0cc0
  X"2f",X"21",X"02",X"00",X"39",X"cd",X"40",X"2f", -- 0cc8
  X"e5",X"3e",X"01",X"cd",X"69",X"2e",X"c1",X"cd", -- 0cd0
  X"4d",X"2f",X"eb",X"21",X"01",X"00",X"cd",X"a8", -- 0cd8
  X"2f",X"7c",X"b5",X"ca",X"14",X"0d",X"21",X"09", -- 0ce0
  X"00",X"e5",X"3e",X"01",X"cd",X"b7",X"26",X"c1", -- 0ce8
  X"21",X"05",X"00",X"39",X"cd",X"4d",X"2f",X"cd", -- 0cf0
  X"40",X"2f",X"e5",X"3e",X"01",X"cd",X"a8",X"24", -- 0cf8
  X"c1",X"21",X"05",X"00",X"39",X"e5",X"cd",X"4d", -- 0d00
  X"2f",X"11",X"01",X"00",X"19",X"d1",X"cd",X"8d", -- 0d08
  X"2f",X"c3",X"a0",X"0d",X"21",X"02",X"00",X"39", -- 0d10
  X"cd",X"40",X"2f",X"e5",X"3e",X"01",X"cd",X"69", -- 0d18
  X"2e",X"c1",X"cd",X"4d",X"2f",X"eb",X"21",X"02", -- 0d20
  X"00",X"cd",X"a8",X"2f",X"7c",X"b5",X"ca",X"5a", -- 0d28
  X"0d",X"21",X"09",X"00",X"e5",X"3e",X"01",X"cd", -- 0d30
  X"b7",X"26",X"c1",X"e1",X"e5",X"cd",X"4d",X"2f", -- 0d38
  X"e5",X"3e",X"01",X"cd",X"e3",X"23",X"c1",X"21", -- 0d40
  X"05",X"00",X"39",X"e5",X"cd",X"4d",X"2f",X"11", -- 0d48
  X"02",X"00",X"19",X"d1",X"cd",X"8d",X"2f",X"c3", -- 0d50
  X"a0",X"0d",X"21",X"02",X"00",X"39",X"cd",X"40", -- 0d58
  X"2f",X"e5",X"3e",X"01",X"cd",X"69",X"2e",X"c1", -- 0d60
  X"cd",X"4d",X"2f",X"7c",X"b5",X"ca",X"92",X"0d", -- 0d68
  X"21",X"09",X"00",X"e5",X"3e",X"01",X"cd",X"b7", -- 0d70
  X"26",X"c1",X"21",X"02",X"00",X"39",X"cd",X"40", -- 0d78
  X"2f",X"e5",X"3e",X"01",X"cd",X"69",X"2e",X"c1", -- 0d80
  X"e5",X"3e",X"01",X"cd",X"68",X"25",X"c1",X"c3", -- 0d88
  X"a0",X"0d",X"af",X"cd",X"d5",X"23",X"21",X"05", -- 0d90
  X"00",X"39",X"cd",X"4d",X"2f",X"33",X"c1",X"c9", -- 0d98
  X"21",X"00",X"00",X"39",X"eb",X"21",X"05",X"00", -- 0da0
  X"39",X"cd",X"4d",X"2f",X"cd",X"8d",X"2f",X"21", -- 0da8
  X"02",X"00",X"39",X"cd",X"40",X"2f",X"e5",X"3e", -- 0db0
  X"01",X"cd",X"7a",X"2e",X"c1",X"cd",X"4d",X"2f", -- 0db8
  X"eb",X"21",X"01",X"00",X"cd",X"a8",X"2f",X"7c", -- 0dc0
  X"b5",X"ca",X"fa",X"0d",X"21",X"2c",X"00",X"e5", -- 0dc8
  X"3e",X"01",X"cd",X"b7",X"26",X"c1",X"21",X"05", -- 0dd0
  X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f", -- 0dd8
  X"e5",X"3e",X"01",X"cd",X"a8",X"24",X"c1",X"21", -- 0de0
  X"05",X"00",X"39",X"e5",X"cd",X"4d",X"2f",X"11", -- 0de8
  X"01",X"00",X"19",X"d1",X"cd",X"8d",X"2f",X"c3", -- 0df0
  X"75",X"0e",X"21",X"02",X"00",X"39",X"cd",X"40", -- 0df8
  X"2f",X"e5",X"3e",X"01",X"cd",X"7a",X"2e",X"c1", -- 0e00
  X"cd",X"4d",X"2f",X"eb",X"21",X"02",X"00",X"cd", -- 0e08
  X"a8",X"2f",X"7c",X"b5",X"ca",X"40",X"0e",X"21", -- 0e10
  X"2c",X"00",X"e5",X"3e",X"01",X"cd",X"b7",X"26", -- 0e18
  X"c1",X"e1",X"e5",X"cd",X"4d",X"2f",X"e5",X"3e", -- 0e20
  X"01",X"cd",X"e3",X"23",X"c1",X"21",X"05",X"00", -- 0e28
  X"39",X"e5",X"cd",X"4d",X"2f",X"11",X"02",X"00", -- 0e30
  X"19",X"d1",X"cd",X"8d",X"2f",X"c3",X"75",X"0e", -- 0e38
  X"21",X"02",X"00",X"39",X"cd",X"40",X"2f",X"e5", -- 0e40
  X"3e",X"01",X"cd",X"7a",X"2e",X"c1",X"cd",X"4d", -- 0e48
  X"2f",X"7c",X"b5",X"ca",X"75",X"0e",X"21",X"2c", -- 0e50
  X"00",X"e5",X"3e",X"01",X"cd",X"b7",X"26",X"c1", -- 0e58
  X"21",X"02",X"00",X"39",X"cd",X"40",X"2f",X"e5", -- 0e60
  X"3e",X"01",X"cd",X"7a",X"2e",X"c1",X"e5",X"3e", -- 0e68
  X"01",X"cd",X"68",X"25",X"c1",X"af",X"cd",X"d5", -- 0e70
  X"23",X"21",X"05",X"00",X"39",X"cd",X"4d",X"2f", -- 0e78
  X"33",X"c1",X"c9",X"21",X"f9",X"0e",X"e5",X"3e", -- 0e80
  X"01",X"cd",X"68",X"25",X"c1",X"21",X"00",X"0f", -- 0e88
  X"e5",X"3e",X"01",X"cd",X"68",X"25",X"c1",X"21", -- 0e90
  X"31",X"0f",X"e5",X"3e",X"01",X"cd",X"68",X"25", -- 0e98
  X"c1",X"af",X"cd",X"d5",X"23",X"21",X"04",X"00", -- 0ea0
  X"39",X"e5",X"21",X"06",X"00",X"39",X"cd",X"4d", -- 0ea8
  X"2f",X"eb",X"21",X"f0",X"ff",X"cd",X"a1",X"2f", -- 0eb0
  X"d1",X"cd",X"8d",X"2f",X"21",X"04",X"00",X"39", -- 0eb8
  X"e5",X"21",X"06",X"00",X"39",X"cd",X"4d",X"2f", -- 0ec0
  X"e5",X"3e",X"01",X"cd",X"37",X"0f",X"c1",X"d1", -- 0ec8
  X"cd",X"8d",X"2f",X"21",X"04",X"00",X"39",X"cd", -- 0ed0
  X"4d",X"2f",X"eb",X"21",X"01",X"00",X"cd",X"04", -- 0ed8
  X"30",X"eb",X"c1",X"e1",X"e5",X"c5",X"cd",X"e5", -- 0ee0
  X"2f",X"7c",X"b5",X"ca",X"f1",X"0e",X"c3",X"bc", -- 0ee8
  X"0e",X"21",X"04",X"00",X"39",X"cd",X"4d",X"2f", -- 0ef0
  X"c9",X"20",X"20",X"20",X"20",X"20",X"20",X"00", -- 0ef8
  X"2b",X"30",X"20",X"2b",X"31",X"20",X"2b",X"32", -- 0f00
  X"20",X"2b",X"33",X"20",X"2b",X"34",X"20",X"2b", -- 0f08
  X"35",X"20",X"2b",X"36",X"20",X"2b",X"37",X"20", -- 0f10
  X"2b",X"38",X"20",X"2b",X"39",X"20",X"2b",X"41", -- 0f18
  X"20",X"2b",X"42",X"20",X"2b",X"43",X"20",X"2b", -- 0f20
  X"44",X"20",X"2b",X"45",X"20",X"2b",X"46",X"20", -- 0f28
  X"00",X"41",X"53",X"43",X"49",X"49",X"00",X"21", -- 0f30
  X"ee",X"ff",X"39",X"f9",X"21",X"20",X"00",X"e5", -- 0f38
  X"3e",X"01",X"cd",X"b7",X"26",X"c1",X"21",X"14", -- 0f40
  X"00",X"39",X"cd",X"4d",X"2f",X"e5",X"3e",X"01", -- 0f48
  X"cd",X"e3",X"23",X"c1",X"21",X"20",X"00",X"e5", -- 0f50
  X"3e",X"01",X"cd",X"b7",X"26",X"c1",X"21",X"00", -- 0f58
  X"00",X"39",X"eb",X"21",X"00",X"00",X"cd",X"8d", -- 0f60
  X"2f",X"d1",X"d5",X"21",X"10",X"00",X"cd",X"c8", -- 0f68
  X"2f",X"7c",X"b5",X"ca",X"aa",X"0f",X"c3",X"8a", -- 0f70
  X"0f",X"21",X"00",X"00",X"39",X"54",X"5d",X"cd", -- 0f78
  X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"c3", -- 0f80
  X"69",X"0f",X"21",X"02",X"00",X"39",X"eb",X"e1", -- 0f88
  X"e5",X"19",X"e5",X"21",X"16",X"00",X"39",X"54", -- 0f90
  X"5d",X"cd",X"4d",X"2f",X"23",X"cd",X"8d",X"2f", -- 0f98
  X"2b",X"cd",X"40",X"2f",X"d1",X"7d",X"12",X"c3", -- 0fa0
  X"79",X"0f",X"21",X"00",X"00",X"39",X"eb",X"21", -- 0fa8
  X"00",X"00",X"cd",X"8d",X"2f",X"d1",X"d5",X"21", -- 0fb0
  X"10",X"00",X"cd",X"c8",X"2f",X"7c",X"b5",X"ca", -- 0fb8
  X"f5",X"0f",X"c3",X"d6",X"0f",X"21",X"00",X"00", -- 0fc0
  X"39",X"54",X"5d",X"cd",X"4d",X"2f",X"23",X"cd", -- 0fc8
  X"8d",X"2f",X"2b",X"c3",X"b5",X"0f",X"21",X"02", -- 0fd0
  X"00",X"39",X"eb",X"e1",X"e5",X"19",X"cd",X"40", -- 0fd8
  X"2f",X"e5",X"3e",X"01",X"cd",X"a8",X"24",X"c1", -- 0fe0
  X"21",X"20",X"00",X"e5",X"3e",X"01",X"cd",X"b7", -- 0fe8
  X"26",X"c1",X"c3",X"c5",X"0f",X"21",X"00",X"00", -- 0ff0
  X"39",X"eb",X"21",X"00",X"00",X"cd",X"8d",X"2f", -- 0ff8
  X"d1",X"d5",X"21",X"10",X"00",X"cd",X"c8",X"2f", -- 1000
  X"7c",X"b5",X"ca",X"5a",X"10",X"c3",X"21",X"10", -- 1008
  X"21",X"00",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 1010
  X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"c3",X"00", -- 1018
  X"10",X"21",X"02",X"00",X"39",X"eb",X"e1",X"e5", -- 1020
  X"19",X"cd",X"40",X"2f",X"e5",X"3e",X"01",X"cd", -- 1028
  X"38",X"1c",X"c1",X"7c",X"b5",X"ca",X"4d",X"10", -- 1030
  X"21",X"02",X"00",X"39",X"eb",X"e1",X"e5",X"19", -- 1038
  X"cd",X"40",X"2f",X"e5",X"3e",X"01",X"cd",X"b7", -- 1040
  X"26",X"c1",X"c3",X"57",X"10",X"21",X"2e",X"00", -- 1048
  X"e5",X"3e",X"01",X"cd",X"b7",X"26",X"c1",X"c3", -- 1050
  X"10",X"10",X"af",X"cd",X"d5",X"23",X"21",X"14", -- 1058
  X"00",X"39",X"cd",X"4d",X"2f",X"eb",X"21",X"12", -- 1060
  X"00",X"39",X"f9",X"eb",X"c9",X"21",X"ae",X"ff", -- 1068
  X"39",X"f9",X"21",X"54",X"00",X"39",X"cd",X"4d", -- 1070
  X"2f",X"cd",X"40",X"2f",X"7c",X"b5",X"ca",X"68", -- 1078
  X"11",X"21",X"54",X"00",X"39",X"cd",X"4d",X"2f", -- 1080
  X"e5",X"21",X"04",X"00",X"39",X"e5",X"21",X"58", -- 1088
  X"00",X"39",X"cd",X"4d",X"2f",X"e5",X"3e",X"03", -- 1090
  X"cd",X"ae",X"1a",X"c1",X"c1",X"c1",X"21",X"00", -- 1098
  X"00",X"39",X"eb",X"21",X"02",X"00",X"39",X"cd", -- 10a0
  X"8d",X"2f",X"e1",X"e5",X"e5",X"3e",X"01",X"cd", -- 10a8
  X"80",X"1d",X"c1",X"7c",X"b5",X"ca",X"d8",X"10", -- 10b0
  X"21",X"56",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 10b8
  X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"e5",X"c1", -- 10c0
  X"e1",X"e5",X"c5",X"e5",X"3e",X"01",X"cd",X"62", -- 10c8
  X"21",X"c1",X"d1",X"7d",X"12",X"c3",X"65",X"11", -- 10d0
  X"e1",X"e5",X"cd",X"40",X"2f",X"eb",X"21",X"27", -- 10d8
  X"00",X"cd",X"a8",X"2f",X"7c",X"b5",X"ca",X"49", -- 10e0
  X"11",X"21",X"00",X"00",X"39",X"54",X"5d",X"cd", -- 10e8
  X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"e1", -- 10f0
  X"e5",X"cd",X"40",X"2f",X"7c",X"b5",X"ca",X"18", -- 10f8
  X"11",X"e1",X"e5",X"cd",X"40",X"2f",X"eb",X"21", -- 1100
  X"27",X"00",X"cd",X"ae",X"2f",X"7c",X"b5",X"ca", -- 1108
  X"18",X"11",X"21",X"01",X"00",X"c3",X"1b",X"11", -- 1110
  X"21",X"00",X"00",X"7c",X"b5",X"ca",X"46",X"11", -- 1118
  X"21",X"56",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 1120
  X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"e5",X"21", -- 1128
  X"02",X"00",X"39",X"54",X"5d",X"cd",X"4d",X"2f", -- 1130
  X"23",X"cd",X"8d",X"2f",X"2b",X"cd",X"40",X"2f", -- 1138
  X"d1",X"7d",X"12",X"c3",X"f7",X"10",X"c3",X"65", -- 1140
  X"11",X"21",X"77",X"11",X"e5",X"3e",X"01",X"cd", -- 1148
  X"68",X"25",X"c1",X"21",X"02",X"00",X"39",X"e5", -- 1150
  X"3e",X"01",X"cd",X"68",X"25",X"c1",X"af",X"cd", -- 1158
  X"d5",X"23",X"c3",X"68",X"11",X"c3",X"72",X"10", -- 1160
  X"21",X"56",X"00",X"39",X"cd",X"4d",X"2f",X"eb", -- 1168
  X"21",X"52",X"00",X"39",X"f9",X"eb",X"c9",X"45", -- 1170
  X"72",X"72",X"6f",X"72",X"2d",X"00",X"c5",X"c5", -- 1178
  X"c5",X"21",X"08",X"00",X"39",X"cd",X"4d",X"2f", -- 1180
  X"cd",X"40",X"2f",X"7c",X"b5",X"c2",X"03",X"12", -- 1188
  X"21",X"c5",X"14",X"e5",X"3e",X"01",X"cd",X"68", -- 1190
  X"25",X"c1",X"af",X"cd",X"d5",X"23",X"21",X"eb", -- 1198
  X"14",X"e5",X"3e",X"01",X"cd",X"68",X"25",X"c1", -- 11a0
  X"af",X"cd",X"d5",X"23",X"21",X"03",X"15",X"e5", -- 11a8
  X"3e",X"01",X"cd",X"68",X"25",X"c1",X"af",X"cd", -- 11b0
  X"d5",X"23",X"21",X"1e",X"15",X"e5",X"3e",X"01", -- 11b8
  X"cd",X"68",X"25",X"c1",X"af",X"cd",X"d5",X"23", -- 11c0
  X"21",X"39",X"15",X"e5",X"3e",X"01",X"cd",X"68", -- 11c8
  X"25",X"c1",X"af",X"cd",X"d5",X"23",X"21",X"55", -- 11d0
  X"15",X"e5",X"3e",X"01",X"cd",X"68",X"25",X"c1", -- 11d8
  X"af",X"cd",X"d5",X"23",X"21",X"74",X"15",X"e5", -- 11e0
  X"3e",X"01",X"cd",X"68",X"25",X"c1",X"af",X"cd", -- 11e8
  X"d5",X"23",X"21",X"90",X"15",X"e5",X"3e",X"01", -- 11f0
  X"cd",X"68",X"25",X"c1",X"af",X"cd",X"d5",X"23", -- 11f8
  X"c3",X"c1",X"14",X"21",X"08",X"00",X"39",X"cd", -- 1200
  X"4d",X"2f",X"cd",X"40",X"2f",X"eb",X"21",X"00", -- 1208
  X"00",X"cd",X"ae",X"2f",X"7c",X"b5",X"ca",X"59", -- 1210
  X"12",X"21",X"08",X"00",X"39",X"cd",X"4d",X"2f", -- 1218
  X"cd",X"40",X"2f",X"e5",X"3e",X"01",X"cd",X"68", -- 1220
  X"1c",X"c1",X"7c",X"b5",X"c2",X"4b",X"12",X"21", -- 1228
  X"08",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40", -- 1230
  X"2f",X"eb",X"21",X"2c",X"00",X"cd",X"a8",X"2f", -- 1238
  X"7c",X"b5",X"c2",X"4b",X"12",X"21",X"00",X"00", -- 1240
  X"c3",X"4e",X"12",X"21",X"01",X"00",X"7c",X"b5", -- 1248
  X"ca",X"59",X"12",X"21",X"01",X"00",X"c3",X"5c", -- 1250
  X"12",X"21",X"00",X"00",X"7c",X"b5",X"ca",X"72", -- 1258
  X"12",X"21",X"08",X"00",X"39",X"54",X"5d",X"cd", -- 1260
  X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"c3", -- 1268
  X"03",X"12",X"21",X"04",X"00",X"39",X"eb",X"21", -- 1270
  X"08",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"8d", -- 1278
  X"2f",X"21",X"04",X"00",X"39",X"cd",X"4d",X"2f", -- 1280
  X"cd",X"40",X"2f",X"eb",X"21",X"00",X"00",X"cd", -- 1288
  X"ae",X"2f",X"7c",X"b5",X"ca",X"cc",X"12",X"21", -- 1290
  X"04",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40", -- 1298
  X"2f",X"e5",X"3e",X"01",X"cd",X"68",X"1c",X"c1", -- 12a0
  X"cd",X"17",X"30",X"7c",X"b5",X"ca",X"cc",X"12", -- 12a8
  X"21",X"04",X"00",X"39",X"cd",X"4d",X"2f",X"cd", -- 12b0
  X"40",X"2f",X"eb",X"21",X"2c",X"00",X"cd",X"ae", -- 12b8
  X"2f",X"7c",X"b5",X"ca",X"cc",X"12",X"21",X"01", -- 12c0
  X"00",X"c3",X"cf",X"12",X"21",X"00",X"00",X"7c", -- 12c8
  X"b5",X"ca",X"e5",X"12",X"21",X"04",X"00",X"39", -- 12d0
  X"54",X"5d",X"cd",X"4d",X"2f",X"23",X"cd",X"8d", -- 12d8
  X"2f",X"2b",X"c3",X"81",X"12",X"21",X"04",X"00", -- 12e0
  X"39",X"cd",X"4d",X"2f",X"eb",X"21",X"00",X"00", -- 12e8
  X"7d",X"12",X"21",X"00",X"00",X"39",X"eb",X"21", -- 12f0
  X"00",X"00",X"cd",X"8d",X"2f",X"21",X"02",X"00", -- 12f8
  X"39",X"eb",X"21",X"00",X"00",X"cd",X"8d",X"2f", -- 1300
  X"c1",X"d1",X"d5",X"c5",X"21",X"ff",X"00",X"cd", -- 1308
  X"bb",X"2f",X"7c",X"b5",X"ca",X"9e",X"14",X"c3", -- 1310
  X"2b",X"13",X"21",X"02",X"00",X"39",X"54",X"5d", -- 1318
  X"cd",X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b", -- 1320
  X"c3",X"08",X"13",X"21",X"08",X"00",X"39",X"cd", -- 1328
  X"4d",X"2f",X"e5",X"21",X"04",X"00",X"39",X"cd", -- 1330
  X"4d",X"2f",X"e5",X"3e",X"01",X"cd",X"58",X"2e", -- 1338
  X"c1",X"e5",X"3e",X"02",X"cd",X"cd",X"1e",X"c1", -- 1340
  X"c1",X"7c",X"b5",X"c2",X"9b",X"14",X"21",X"b0", -- 1348
  X"15",X"e5",X"3e",X"01",X"cd",X"68",X"25",X"c1", -- 1350
  X"c1",X"e1",X"e5",X"c5",X"e5",X"3e",X"01",X"cd", -- 1358
  X"58",X"2e",X"c1",X"e5",X"3e",X"01",X"cd",X"68", -- 1360
  X"25",X"c1",X"c1",X"e1",X"e5",X"c5",X"e5",X"3e", -- 1368
  X"01",X"cd",X"69",X"2e",X"c1",X"cd",X"4d",X"2f", -- 1370
  X"eb",X"21",X"01",X"00",X"cd",X"a8",X"2f",X"7c", -- 1378
  X"b5",X"ca",X"9b",X"13",X"21",X"09",X"00",X"e5", -- 1380
  X"3e",X"01",X"cd",X"b7",X"26",X"c1",X"21",X"b7", -- 1388
  X"15",X"e5",X"3e",X"01",X"cd",X"68",X"25",X"c1", -- 1390
  X"c3",X"fb",X"13",X"c1",X"e1",X"e5",X"c5",X"e5", -- 1398
  X"3e",X"01",X"cd",X"69",X"2e",X"c1",X"cd",X"4d", -- 13a0
  X"2f",X"eb",X"21",X"02",X"00",X"cd",X"a8",X"2f", -- 13a8
  X"7c",X"b5",X"ca",X"cc",X"13",X"21",X"09",X"00", -- 13b0
  X"e5",X"3e",X"01",X"cd",X"b7",X"26",X"c1",X"21", -- 13b8
  X"ba",X"15",X"e5",X"3e",X"01",X"cd",X"68",X"25", -- 13c0
  X"c1",X"c3",X"fb",X"13",X"c1",X"e1",X"e5",X"c5", -- 13c8
  X"e5",X"3e",X"01",X"cd",X"69",X"2e",X"c1",X"cd", -- 13d0
  X"4d",X"2f",X"7c",X"b5",X"ca",X"fb",X"13",X"21", -- 13d8
  X"09",X"00",X"e5",X"3e",X"01",X"cd",X"b7",X"26", -- 13e0
  X"c1",X"c1",X"e1",X"e5",X"c5",X"e5",X"3e",X"01", -- 13e8
  X"cd",X"69",X"2e",X"c1",X"e5",X"3e",X"01",X"cd", -- 13f0
  X"68",X"25",X"c1",X"c1",X"e1",X"e5",X"c5",X"e5", -- 13f8
  X"3e",X"01",X"cd",X"7a",X"2e",X"c1",X"cd",X"4d", -- 1400
  X"2f",X"eb",X"21",X"01",X"00",X"cd",X"a8",X"2f", -- 1408
  X"7c",X"b5",X"ca",X"2c",X"14",X"21",X"2c",X"00", -- 1410
  X"e5",X"3e",X"01",X"cd",X"b7",X"26",X"c1",X"21", -- 1418
  X"bf",X"15",X"e5",X"3e",X"01",X"cd",X"68",X"25", -- 1420
  X"c1",X"c3",X"8c",X"14",X"c1",X"e1",X"e5",X"c5", -- 1428
  X"e5",X"3e",X"01",X"cd",X"7a",X"2e",X"c1",X"cd", -- 1430
  X"4d",X"2f",X"eb",X"21",X"02",X"00",X"cd",X"a8", -- 1438
  X"2f",X"7c",X"b5",X"ca",X"5d",X"14",X"21",X"2c", -- 1440
  X"00",X"e5",X"3e",X"01",X"cd",X"b7",X"26",X"c1", -- 1448
  X"21",X"c2",X"15",X"e5",X"3e",X"01",X"cd",X"68", -- 1450
  X"25",X"c1",X"c3",X"8c",X"14",X"c1",X"e1",X"e5", -- 1458
  X"c5",X"e5",X"3e",X"01",X"cd",X"7a",X"2e",X"c1", -- 1460
  X"cd",X"4d",X"2f",X"7c",X"b5",X"ca",X"8c",X"14", -- 1468
  X"21",X"2c",X"00",X"e5",X"3e",X"01",X"cd",X"b7", -- 1470
  X"26",X"c1",X"c1",X"e1",X"e5",X"c5",X"e5",X"3e", -- 1478
  X"01",X"cd",X"7a",X"2e",X"c1",X"e5",X"3e",X"01", -- 1480
  X"cd",X"68",X"25",X"c1",X"af",X"cd",X"d5",X"23", -- 1488
  X"21",X"00",X"00",X"39",X"eb",X"21",X"01",X"00", -- 1490
  X"cd",X"8d",X"2f",X"c3",X"1a",X"13",X"e1",X"e5", -- 1498
  X"7c",X"b5",X"c2",X"c1",X"14",X"21",X"c7",X"15", -- 14a0
  X"e5",X"3e",X"01",X"cd",X"68",X"25",X"c1",X"21", -- 14a8
  X"08",X"00",X"39",X"cd",X"4d",X"2f",X"e5",X"3e", -- 14b0
  X"01",X"cd",X"68",X"25",X"c1",X"af",X"cd",X"d5", -- 14b8
  X"23",X"c1",X"c1",X"c1",X"c9",X"20",X"20",X"20", -- 14c0
  X"20",X"20",X"20",X"78",X"78",X"78",X"78",X"20", -- 14c8
  X"20",X"20",X"20",X"20",X"43",X"68",X"61",X"6e", -- 14d0
  X"67",X"65",X"20",X"63",X"75",X"72",X"72",X"65", -- 14d8
  X"6e",X"74",X"20",X"61",X"64",X"64",X"72",X"65", -- 14e0
  X"73",X"73",X"00",X"20",X"20",X"20",X"20",X"20", -- 14e8
  X"20",X"6d",X"6e",X"65",X"6d",X"6f",X"6e",X"69", -- 14f0
  X"63",X"20",X"41",X"73",X"73",X"65",X"6d",X"62", -- 14f8
  X"6c",X"65",X"00",X"20",X"20",X"20",X"20",X"20", -- 1500
  X"20",X"4c",X"49",X"53",X"54",X"20",X"20",X"20", -- 1508
  X"20",X"20",X"44",X"69",X"73",X"61",X"73",X"73", -- 1510
  X"65",X"6d",X"62",X"6c",X"65",X"00",X"20",X"20", -- 1518
  X"20",X"20",X"20",X"20",X"44",X"45",X"46",X"49", -- 1520
  X"4e",X"45",X"20",X"20",X"20",X"44",X"65",X"66", -- 1528
  X"69",X"6e",X"65",X"20",X"64",X"61",X"74",X"61", -- 1530
  X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"44", -- 1538
  X"55",X"4d",X"50",X"20",X"20",X"20",X"20",X"20", -- 1540
  X"44",X"69",X"73",X"70",X"6c",X"61",X"79",X"20", -- 1548
  X"64",X"61",X"74",X"61",X"00",X"20",X"20",X"20", -- 1550
  X"20",X"20",X"20",X"45",X"58",X"45",X"43",X"20", -- 1558
  X"20",X"20",X"20",X"20",X"45",X"78",X"65",X"63", -- 1560
  X"75",X"74",X"65",X"20",X"70",X"72",X"6f",X"67", -- 1568
  X"72",X"61",X"6d",X"00",X"20",X"20",X"20",X"20", -- 1570
  X"20",X"20",X"48",X"45",X"4c",X"50",X"20",X"20", -- 1578
  X"20",X"20",X"20",X"44",X"69",X"73",X"70",X"6c", -- 1580
  X"61",X"79",X"20",X"68",X"65",X"6c",X"70",X"00", -- 1588
  X"20",X"20",X"20",X"20",X"20",X"20",X"53",X"59", -- 1590
  X"53",X"54",X"45",X"4d",X"20",X"20",X"20",X"52", -- 1598
  X"65",X"74",X"75",X"72",X"6e",X"20",X"74",X"6f", -- 15a0
  X"20",X"73",X"79",X"73",X"74",X"65",X"6d",X"00", -- 15a8
  X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"78", -- 15b0
  X"78",X"00",X"78",X"78",X"78",X"78",X"00",X"78", -- 15b8
  X"78",X"00",X"78",X"78",X"78",X"78",X"00",X"45", -- 15c0
  X"52",X"52",X"4f",X"52",X"2d",X"00",X"3b",X"c5", -- 15c8
  X"c5",X"21",X"04",X"00",X"39",X"eb",X"21",X"ff", -- 15d0
  X"00",X"7d",X"12",X"21",X"00",X"00",X"39",X"eb", -- 15d8
  X"21",X"00",X"00",X"cd",X"8d",X"2f",X"21",X"04", -- 15e0
  X"00",X"39",X"54",X"5d",X"cd",X"40",X"2f",X"2b", -- 15e8
  X"7d",X"12",X"23",X"7c",X"b5",X"ca",X"0b",X"16", -- 15f0
  X"d1",X"d5",X"21",X"00",X"00",X"cd",X"a8",X"2f", -- 15f8
  X"7c",X"b5",X"ca",X"0b",X"16",X"21",X"01",X"00", -- 1600
  X"c3",X"0e",X"16",X"21",X"00",X"00",X"7c",X"b5", -- 1608
  X"ca",X"30",X"17",X"21",X"0b",X"00",X"39",X"cd", -- 1610
  X"4d",X"2f",X"e5",X"21",X"06",X"00",X"39",X"cd", -- 1618
  X"40",X"2f",X"e5",X"3e",X"01",X"cd",X"58",X"2e", -- 1620
  X"c1",X"e5",X"3e",X"02",X"cd",X"cd",X"1e",X"c1", -- 1628
  X"c1",X"7c",X"b5",X"c2",X"2d",X"17",X"21",X"09", -- 1630
  X"00",X"39",X"cd",X"4d",X"2f",X"e5",X"21",X"06", -- 1638
  X"00",X"39",X"cd",X"40",X"2f",X"e5",X"3e",X"01", -- 1640
  X"cd",X"69",X"2e",X"c1",X"e5",X"3e",X"02",X"cd", -- 1648
  X"cd",X"1e",X"c1",X"c1",X"eb",X"21",X"00",X"00", -- 1650
  X"cd",X"a8",X"2f",X"7c",X"b5",X"c2",X"a4",X"16", -- 1658
  X"21",X"09",X"00",X"39",X"cd",X"4d",X"2f",X"e5", -- 1660
  X"3e",X"01",X"cd",X"80",X"1d",X"c1",X"7c",X"b5", -- 1668
  X"ca",X"96",X"16",X"21",X"04",X"00",X"39",X"cd", -- 1670
  X"40",X"2f",X"e5",X"3e",X"01",X"cd",X"69",X"2e", -- 1678
  X"c1",X"cd",X"4d",X"2f",X"eb",X"21",X"02",X"00", -- 1680
  X"cd",X"bb",X"2f",X"7c",X"b5",X"ca",X"96",X"16", -- 1688
  X"21",X"01",X"00",X"c3",X"99",X"16",X"21",X"00", -- 1690
  X"00",X"7c",X"b5",X"c2",X"a4",X"16",X"21",X"00", -- 1698
  X"00",X"c3",X"a7",X"16",X"21",X"01",X"00",X"7c", -- 16a0
  X"b5",X"ca",X"2d",X"17",X"21",X"07",X"00",X"39", -- 16a8
  X"cd",X"4d",X"2f",X"e5",X"21",X"06",X"00",X"39", -- 16b0
  X"cd",X"40",X"2f",X"e5",X"3e",X"01",X"cd",X"7a", -- 16b8
  X"2e",X"c1",X"e5",X"3e",X"02",X"cd",X"cd",X"1e", -- 16c0
  X"c1",X"c1",X"eb",X"21",X"00",X"00",X"cd",X"a8", -- 16c8
  X"2f",X"7c",X"b5",X"c2",X"1a",X"17",X"21",X"07", -- 16d0
  X"00",X"39",X"cd",X"4d",X"2f",X"e5",X"3e",X"01", -- 16d8
  X"cd",X"80",X"1d",X"c1",X"7c",X"b5",X"ca",X"0c", -- 16e0
  X"17",X"21",X"04",X"00",X"39",X"cd",X"40",X"2f", -- 16e8
  X"e5",X"3e",X"01",X"cd",X"7a",X"2e",X"c1",X"cd", -- 16f0
  X"4d",X"2f",X"eb",X"21",X"02",X"00",X"cd",X"bb", -- 16f8
  X"2f",X"7c",X"b5",X"ca",X"0c",X"17",X"21",X"01", -- 1700
  X"00",X"c3",X"0f",X"17",X"21",X"00",X"00",X"7c", -- 1708
  X"b5",X"c2",X"1a",X"17",X"21",X"00",X"00",X"c3", -- 1710
  X"1d",X"17",X"21",X"01",X"00",X"7c",X"b5",X"ca", -- 1718
  X"2d",X"17",X"21",X"00",X"00",X"39",X"eb",X"21", -- 1720
  X"01",X"00",X"cd",X"8d",X"2f",X"c3",X"e6",X"15", -- 1728
  X"e1",X"e5",X"7c",X"b5",X"c2",X"ac",X"17",X"21", -- 1730
  X"08",X"19",X"e5",X"3e",X"01",X"cd",X"68",X"25", -- 1738
  X"c1",X"21",X"0b",X"00",X"39",X"cd",X"4d",X"2f", -- 1740
  X"e5",X"3e",X"01",X"cd",X"68",X"25",X"c1",X"21", -- 1748
  X"20",X"00",X"e5",X"3e",X"01",X"cd",X"b7",X"26", -- 1750
  X"c1",X"21",X"09",X"00",X"39",X"cd",X"4d",X"2f", -- 1758
  X"cd",X"40",X"2f",X"7c",X"b5",X"ca",X"76",X"17", -- 1760
  X"21",X"09",X"00",X"39",X"cd",X"4d",X"2f",X"e5", -- 1768
  X"3e",X"01",X"cd",X"68",X"25",X"c1",X"21",X"07", -- 1770
  X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f", -- 1778
  X"7c",X"b5",X"ca",X"9d",X"17",X"21",X"2c",X"00", -- 1780
  X"e5",X"3e",X"01",X"cd",X"b7",X"26",X"c1",X"21", -- 1788
  X"07",X"00",X"39",X"cd",X"4d",X"2f",X"e5",X"3e", -- 1790
  X"01",X"cd",X"68",X"25",X"c1",X"af",X"cd",X"d5", -- 1798
  X"23",X"21",X"0d",X"00",X"39",X"cd",X"4d",X"2f", -- 17a0
  X"33",X"c1",X"c1",X"c9",X"21",X"04",X"00",X"39", -- 17a8
  X"54",X"5d",X"cd",X"40",X"2f",X"23",X"7d",X"12", -- 17b0
  X"2b",X"21",X"0d",X"00",X"39",X"54",X"5d",X"cd", -- 17b8
  X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"eb", -- 17c0
  X"21",X"04",X"00",X"39",X"cd",X"40",X"2f",X"7d", -- 17c8
  X"12",X"21",X"02",X"00",X"39",X"eb",X"21",X"0d", -- 17d0
  X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"8d",X"2f", -- 17d8
  X"21",X"04",X"00",X"39",X"cd",X"40",X"2f",X"e5", -- 17e0
  X"3e",X"01",X"cd",X"69",X"2e",X"c1",X"cd",X"4d", -- 17e8
  X"2f",X"eb",X"21",X"01",X"00",X"cd",X"a8",X"2f", -- 17f0
  X"7c",X"b5",X"ca",X"29",X"18",X"21",X"0d",X"00", -- 17f8
  X"39",X"cd",X"4d",X"2f",X"e5",X"21",X"0b",X"00", -- 1800
  X"39",X"cd",X"4d",X"2f",X"e5",X"3e",X"01",X"cd", -- 1808
  X"62",X"21",X"c1",X"d1",X"7d",X"12",X"21",X"0d", -- 1810
  X"00",X"39",X"e5",X"cd",X"4d",X"2f",X"11",X"01", -- 1818
  X"00",X"19",X"d1",X"cd",X"8d",X"2f",X"c3",X"fd", -- 1820
  X"18",X"21",X"04",X"00",X"39",X"cd",X"40",X"2f", -- 1828
  X"e5",X"3e",X"01",X"cd",X"7a",X"2e",X"c1",X"cd", -- 1830
  X"4d",X"2f",X"eb",X"21",X"01",X"00",X"cd",X"a8", -- 1838
  X"2f",X"7c",X"b5",X"ca",X"72",X"18",X"21",X"0d", -- 1840
  X"00",X"39",X"cd",X"4d",X"2f",X"e5",X"21",X"09", -- 1848
  X"00",X"39",X"cd",X"4d",X"2f",X"e5",X"3e",X"01", -- 1850
  X"cd",X"62",X"21",X"c1",X"d1",X"7d",X"12",X"21", -- 1858
  X"0d",X"00",X"39",X"e5",X"cd",X"4d",X"2f",X"11", -- 1860
  X"01",X"00",X"19",X"d1",X"cd",X"8d",X"2f",X"c3", -- 1868
  X"fd",X"18",X"21",X"04",X"00",X"39",X"cd",X"40", -- 1870
  X"2f",X"e5",X"3e",X"01",X"cd",X"69",X"2e",X"c1", -- 1878
  X"cd",X"4d",X"2f",X"eb",X"21",X"02",X"00",X"cd", -- 1880
  X"a8",X"2f",X"7c",X"b5",X"ca",X"b9",X"18",X"c1", -- 1888
  X"e1",X"e5",X"c5",X"e5",X"21",X"0b",X"00",X"39", -- 1890
  X"cd",X"4d",X"2f",X"e5",X"3e",X"01",X"cd",X"9b", -- 1898
  X"22",X"c1",X"d1",X"cd",X"8d",X"2f",X"21",X"0d", -- 18a0
  X"00",X"39",X"e5",X"cd",X"4d",X"2f",X"11",X"02", -- 18a8
  X"00",X"19",X"d1",X"cd",X"8d",X"2f",X"c3",X"fd", -- 18b0
  X"18",X"21",X"04",X"00",X"39",X"cd",X"40",X"2f", -- 18b8
  X"e5",X"3e",X"01",X"cd",X"7a",X"2e",X"c1",X"cd", -- 18c0
  X"4d",X"2f",X"eb",X"21",X"02",X"00",X"cd",X"a8", -- 18c8
  X"2f",X"7c",X"b5",X"ca",X"fd",X"18",X"c1",X"e1", -- 18d0
  X"e5",X"c5",X"e5",X"21",X"09",X"00",X"39",X"cd", -- 18d8
  X"4d",X"2f",X"e5",X"3e",X"01",X"cd",X"9b",X"22", -- 18e0
  X"c1",X"d1",X"cd",X"8d",X"2f",X"21",X"0d",X"00", -- 18e8
  X"39",X"e5",X"cd",X"4d",X"2f",X"11",X"02",X"00", -- 18f0
  X"19",X"d1",X"cd",X"8d",X"2f",X"21",X"0d",X"00", -- 18f8
  X"39",X"cd",X"4d",X"2f",X"33",X"c1",X"c1",X"c9", -- 1900
  X"45",X"52",X"52",X"4f",X"52",X"2d",X"00",X"21", -- 1908
  X"5b",X"00",X"e5",X"3e",X"01",X"cd",X"b7",X"26", -- 1910
  X"c1",X"c1",X"e1",X"e5",X"c5",X"e5",X"3e",X"01", -- 1918
  X"cd",X"e3",X"23",X"c1",X"21",X"5d",X"00",X"e5", -- 1920
  X"3e",X"01",X"cd",X"b7",X"26",X"c1",X"c9",X"21", -- 1928
  X"06",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40", -- 1930
  X"2f",X"eb",X"21",X"00",X"00",X"cd",X"ae",X"2f", -- 1938
  X"7c",X"b5",X"ca",X"85",X"19",X"21",X"06",X"00", -- 1940
  X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"e5", -- 1948
  X"3e",X"01",X"cd",X"68",X"1c",X"c1",X"7c",X"b5", -- 1950
  X"c2",X"77",X"19",X"21",X"06",X"00",X"39",X"cd", -- 1958
  X"4d",X"2f",X"cd",X"40",X"2f",X"eb",X"21",X"2c", -- 1960
  X"00",X"cd",X"a8",X"2f",X"7c",X"b5",X"c2",X"77", -- 1968
  X"19",X"21",X"00",X"00",X"c3",X"7a",X"19",X"21", -- 1970
  X"01",X"00",X"7c",X"b5",X"ca",X"85",X"19",X"21", -- 1978
  X"01",X"00",X"c3",X"88",X"19",X"21",X"00",X"00", -- 1980
  X"7c",X"b5",X"ca",X"9e",X"19",X"21",X"06",X"00", -- 1988
  X"39",X"54",X"5d",X"cd",X"4d",X"2f",X"23",X"cd", -- 1990
  X"8d",X"2f",X"2b",X"c3",X"2f",X"19",X"21",X"06", -- 1998
  X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f", -- 19a0
  X"eb",X"21",X"00",X"00",X"cd",X"ae",X"2f",X"7c", -- 19a8
  X"b5",X"ca",X"e9",X"19",X"21",X"06",X"00",X"39", -- 19b0
  X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"e5",X"3e", -- 19b8
  X"01",X"cd",X"68",X"1c",X"c1",X"cd",X"17",X"30", -- 19c0
  X"7c",X"b5",X"ca",X"e9",X"19",X"21",X"06",X"00", -- 19c8
  X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"eb", -- 19d0
  X"21",X"2c",X"00",X"cd",X"ae",X"2f",X"7c",X"b5", -- 19d8
  X"ca",X"e9",X"19",X"21",X"01",X"00",X"c3",X"ec", -- 19e0
  X"19",X"21",X"00",X"00",X"7c",X"b5",X"ca",X"17", -- 19e8
  X"1a",X"21",X"04",X"00",X"39",X"54",X"5d",X"cd", -- 19f0
  X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"e5", -- 19f8
  X"21",X"08",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 1a00
  X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"cd",X"40", -- 1a08
  X"2f",X"d1",X"7d",X"12",X"c3",X"9e",X"19",X"21", -- 1a10
  X"04",X"00",X"39",X"cd",X"4d",X"2f",X"eb",X"21", -- 1a18
  X"00",X"00",X"7d",X"12",X"21",X"06",X"00",X"39", -- 1a20
  X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"eb",X"21", -- 1a28
  X"00",X"00",X"cd",X"ae",X"2f",X"7c",X"b5",X"ca", -- 1a30
  X"56",X"1a",X"21",X"06",X"00",X"39",X"cd",X"4d", -- 1a38
  X"2f",X"cd",X"40",X"2f",X"eb",X"21",X"20",X"00", -- 1a40
  X"cd",X"a8",X"2f",X"7c",X"b5",X"ca",X"56",X"1a", -- 1a48
  X"21",X"01",X"00",X"c3",X"59",X"1a",X"21",X"00", -- 1a50
  X"00",X"7c",X"b5",X"ca",X"6f",X"1a",X"21",X"06", -- 1a58
  X"00",X"39",X"54",X"5d",X"cd",X"4d",X"2f",X"23", -- 1a60
  X"cd",X"8d",X"2f",X"2b",X"c3",X"24",X"1a",X"21", -- 1a68
  X"06",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40", -- 1a70
  X"2f",X"7c",X"b5",X"ca",X"a4",X"1a",X"21",X"02", -- 1a78
  X"00",X"39",X"54",X"5d",X"cd",X"4d",X"2f",X"23", -- 1a80
  X"cd",X"8d",X"2f",X"2b",X"e5",X"21",X"08",X"00", -- 1a88
  X"39",X"54",X"5d",X"cd",X"4d",X"2f",X"23",X"cd", -- 1a90
  X"8d",X"2f",X"2b",X"cd",X"40",X"2f",X"d1",X"7d", -- 1a98
  X"12",X"c3",X"6f",X"1a",X"c1",X"d1",X"d5",X"c5", -- 1aa0
  X"21",X"00",X"00",X"7d",X"12",X"c9",X"21",X"06", -- 1aa8
  X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f", -- 1ab0
  X"eb",X"21",X"00",X"00",X"cd",X"ae",X"2f",X"7c", -- 1ab8
  X"b5",X"ca",X"e0",X"1a",X"21",X"06",X"00",X"39", -- 1ac0
  X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"eb",X"21", -- 1ac8
  X"20",X"00",X"cd",X"a8",X"2f",X"7c",X"b5",X"ca", -- 1ad0
  X"e0",X"1a",X"21",X"01",X"00",X"c3",X"e3",X"1a", -- 1ad8
  X"21",X"00",X"00",X"7c",X"b5",X"ca",X"f9",X"1a", -- 1ae0
  X"21",X"06",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 1ae8
  X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"c3",X"ae", -- 1af0
  X"1a",X"21",X"06",X"00",X"39",X"cd",X"4d",X"2f", -- 1af8
  X"cd",X"40",X"2f",X"eb",X"21",X"00",X"00",X"cd", -- 1b00
  X"ae",X"2f",X"7c",X"b5",X"ca",X"2b",X"1b",X"21", -- 1b08
  X"06",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40", -- 1b10
  X"2f",X"eb",X"21",X"2c",X"00",X"cd",X"ae",X"2f", -- 1b18
  X"7c",X"b5",X"ca",X"2b",X"1b",X"21",X"01",X"00", -- 1b20
  X"c3",X"2e",X"1b",X"21",X"00",X"00",X"7c",X"b5", -- 1b28
  X"ca",X"59",X"1b",X"21",X"04",X"00",X"39",X"54", -- 1b30
  X"5d",X"cd",X"4d",X"2f",X"23",X"cd",X"8d",X"2f", -- 1b38
  X"2b",X"e5",X"21",X"08",X"00",X"39",X"54",X"5d", -- 1b40
  X"cd",X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b", -- 1b48
  X"cd",X"40",X"2f",X"d1",X"7d",X"12",X"c3",X"f9", -- 1b50
  X"1a",X"21",X"04",X"00",X"39",X"cd",X"4d",X"2f", -- 1b58
  X"eb",X"21",X"00",X"00",X"7d",X"12",X"21",X"06", -- 1b60
  X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f", -- 1b68
  X"eb",X"21",X"00",X"00",X"cd",X"ae",X"2f",X"7c", -- 1b70
  X"b5",X"ca",X"98",X"1b",X"21",X"06",X"00",X"39", -- 1b78
  X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"eb",X"21", -- 1b80
  X"2c",X"00",X"cd",X"a8",X"2f",X"7c",X"b5",X"ca", -- 1b88
  X"98",X"1b",X"21",X"01",X"00",X"c3",X"9b",X"1b", -- 1b90
  X"21",X"00",X"00",X"7c",X"b5",X"ca",X"ae",X"1b", -- 1b98
  X"21",X"06",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 1ba0
  X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"21",X"06", -- 1ba8
  X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f", -- 1bb0
  X"eb",X"21",X"00",X"00",X"cd",X"ae",X"2f",X"7c", -- 1bb8
  X"b5",X"ca",X"e0",X"1b",X"21",X"06",X"00",X"39", -- 1bc0
  X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"eb",X"21", -- 1bc8
  X"20",X"00",X"cd",X"a8",X"2f",X"7c",X"b5",X"ca", -- 1bd0
  X"e0",X"1b",X"21",X"01",X"00",X"c3",X"e3",X"1b", -- 1bd8
  X"21",X"00",X"00",X"7c",X"b5",X"ca",X"f9",X"1b", -- 1be0
  X"21",X"06",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 1be8
  X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"c3",X"ae", -- 1bf0
  X"1b",X"21",X"06",X"00",X"39",X"cd",X"4d",X"2f", -- 1bf8
  X"cd",X"40",X"2f",X"7c",X"b5",X"ca",X"2e",X"1c", -- 1c00
  X"21",X"02",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 1c08
  X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"e5",X"21", -- 1c10
  X"08",X"00",X"39",X"54",X"5d",X"cd",X"4d",X"2f", -- 1c18
  X"23",X"cd",X"8d",X"2f",X"2b",X"cd",X"40",X"2f", -- 1c20
  X"d1",X"7d",X"12",X"c3",X"f9",X"1b",X"c1",X"d1", -- 1c28
  X"d5",X"c5",X"21",X"00",X"00",X"7d",X"12",X"c9", -- 1c30
  X"21",X"02",X"00",X"39",X"cd",X"40",X"2f",X"eb", -- 1c38
  X"21",X"20",X"00",X"cd",X"c2",X"2f",X"7c",X"b5", -- 1c40
  X"ca",X"64",X"1c",X"21",X"02",X"00",X"39",X"cd", -- 1c48
  X"40",X"2f",X"eb",X"21",X"7e",X"00",X"cd",X"bb", -- 1c50
  X"2f",X"7c",X"b5",X"ca",X"64",X"1c",X"21",X"01", -- 1c58
  X"00",X"c3",X"67",X"1c",X"21",X"00",X"00",X"c9", -- 1c60
  X"21",X"02",X"00",X"39",X"cd",X"40",X"2f",X"eb", -- 1c68
  X"21",X"20",X"00",X"cd",X"bb",X"2f",X"7c",X"b5", -- 1c70
  X"ca",X"d6",X"1c",X"21",X"02",X"00",X"39",X"cd", -- 1c78
  X"40",X"2f",X"eb",X"21",X"20",X"00",X"cd",X"a8", -- 1c80
  X"2f",X"7c",X"b5",X"c2",X"c8",X"1c",X"21",X"02", -- 1c88
  X"00",X"39",X"cd",X"40",X"2f",X"eb",X"21",X"0d", -- 1c90
  X"00",X"cd",X"bb",X"2f",X"7c",X"b5",X"ca",X"ba", -- 1c98
  X"1c",X"21",X"02",X"00",X"39",X"cd",X"40",X"2f", -- 1ca0
  X"eb",X"21",X"09",X"00",X"cd",X"c2",X"2f",X"7c", -- 1ca8
  X"b5",X"ca",X"ba",X"1c",X"21",X"01",X"00",X"c3", -- 1cb0
  X"bd",X"1c",X"21",X"00",X"00",X"7c",X"b5",X"c2", -- 1cb8
  X"c8",X"1c",X"21",X"00",X"00",X"c3",X"cb",X"1c", -- 1cc0
  X"21",X"01",X"00",X"7c",X"b5",X"ca",X"d6",X"1c", -- 1cc8
  X"21",X"01",X"00",X"c3",X"d9",X"1c",X"21",X"00", -- 1cd0
  X"00",X"c9",X"21",X"02",X"00",X"39",X"cd",X"40", -- 1cd8
  X"2f",X"eb",X"21",X"66",X"00",X"cd",X"bb",X"2f", -- 1ce0
  X"7c",X"b5",X"ca",X"06",X"1d",X"21",X"02",X"00", -- 1ce8
  X"39",X"cd",X"40",X"2f",X"eb",X"21",X"61",X"00", -- 1cf0
  X"cd",X"c2",X"2f",X"7c",X"b5",X"ca",X"06",X"1d", -- 1cf8
  X"21",X"01",X"00",X"c3",X"09",X"1d",X"21",X"00", -- 1d00
  X"00",X"7c",X"b5",X"c2",X"7c",X"1d",X"21",X"02", -- 1d08
  X"00",X"39",X"cd",X"40",X"2f",X"eb",X"21",X"46", -- 1d10
  X"00",X"cd",X"bb",X"2f",X"7c",X"b5",X"ca",X"3a", -- 1d18
  X"1d",X"21",X"02",X"00",X"39",X"cd",X"40",X"2f", -- 1d20
  X"eb",X"21",X"41",X"00",X"cd",X"c2",X"2f",X"7c", -- 1d28
  X"b5",X"ca",X"3a",X"1d",X"21",X"01",X"00",X"c3", -- 1d30
  X"3d",X"1d",X"21",X"00",X"00",X"7c",X"b5",X"c2", -- 1d38
  X"7c",X"1d",X"21",X"02",X"00",X"39",X"cd",X"40", -- 1d40
  X"2f",X"eb",X"21",X"39",X"00",X"cd",X"bb",X"2f", -- 1d48
  X"7c",X"b5",X"ca",X"6e",X"1d",X"21",X"02",X"00", -- 1d50
  X"39",X"cd",X"40",X"2f",X"eb",X"21",X"30",X"00", -- 1d58
  X"cd",X"c2",X"2f",X"7c",X"b5",X"ca",X"6e",X"1d", -- 1d60
  X"21",X"01",X"00",X"c3",X"71",X"1d",X"21",X"00", -- 1d68
  X"00",X"7c",X"b5",X"c2",X"7c",X"1d",X"21",X"00", -- 1d70
  X"00",X"c3",X"7f",X"1d",X"21",X"01",X"00",X"c9", -- 1d78
  X"c1",X"e1",X"e5",X"c5",X"cd",X"40",X"2f",X"eb", -- 1d80
  X"21",X"00",X"00",X"cd",X"a8",X"2f",X"7c",X"b5", -- 1d88
  X"c2",X"b5",X"1d",X"c1",X"e1",X"e5",X"c5",X"e5", -- 1d90
  X"21",X"8e",X"1e",X"e5",X"3e",X"02",X"cd",X"cd", -- 1d98
  X"1e",X"c1",X"c1",X"eb",X"21",X"00",X"00",X"cd", -- 1da0
  X"a8",X"2f",X"7c",X"b5",X"c2",X"b5",X"1d",X"21", -- 1da8
  X"00",X"00",X"c3",X"b8",X"1d",X"21",X"01",X"00", -- 1db0
  X"7c",X"b5",X"ca",X"c1",X"1d",X"21",X"00",X"00", -- 1db8
  X"c9",X"c1",X"e1",X"e5",X"c5",X"e5",X"21",X"92", -- 1dc0
  X"1e",X"e5",X"3e",X"02",X"cd",X"cd",X"1e",X"c1", -- 1dc8
  X"c1",X"eb",X"21",X"00",X"00",X"cd",X"a8",X"2f", -- 1dd0
  X"7c",X"b5",X"c2",X"ff",X"1d",X"c1",X"e1",X"e5", -- 1dd8
  X"c5",X"e5",X"21",X"96",X"1e",X"e5",X"3e",X"02", -- 1de0
  X"cd",X"cd",X"1e",X"c1",X"c1",X"eb",X"21",X"00", -- 1de8
  X"00",X"cd",X"a8",X"2f",X"7c",X"b5",X"c2",X"ff", -- 1df0
  X"1d",X"21",X"00",X"00",X"c3",X"02",X"1e",X"21", -- 1df8
  X"01",X"00",X"7c",X"b5",X"ca",X"0b",X"1e",X"21", -- 1e00
  X"00",X"00",X"c9",X"c1",X"e1",X"e5",X"c5",X"e5", -- 1e08
  X"21",X"99",X"1e",X"e5",X"3e",X"02",X"cd",X"cd", -- 1e10
  X"1e",X"c1",X"c1",X"eb",X"21",X"00",X"00",X"cd", -- 1e18
  X"a8",X"2f",X"7c",X"b5",X"c2",X"49",X"1e",X"c1", -- 1e20
  X"e1",X"e5",X"c5",X"e5",X"21",X"9d",X"1e",X"e5", -- 1e28
  X"3e",X"02",X"cd",X"cd",X"1e",X"c1",X"c1",X"eb", -- 1e30
  X"21",X"00",X"00",X"cd",X"a8",X"2f",X"7c",X"b5", -- 1e38
  X"c2",X"49",X"1e",X"21",X"00",X"00",X"c3",X"4c", -- 1e40
  X"1e",X"21",X"01",X"00",X"7c",X"b5",X"ca",X"55", -- 1e48
  X"1e",X"21",X"00",X"00",X"c9",X"c1",X"e1",X"e5", -- 1e50
  X"c5",X"cd",X"40",X"2f",X"e5",X"3e",X"01",X"cd", -- 1e58
  X"da",X"1c",X"c1",X"7c",X"b5",X"ca",X"79",X"1e", -- 1e60
  X"21",X"02",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 1e68
  X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"c3",X"55", -- 1e70
  X"1e",X"c1",X"e1",X"e5",X"c5",X"cd",X"40",X"2f", -- 1e78
  X"7c",X"b5",X"c2",X"89",X"1e",X"21",X"01",X"00", -- 1e80
  X"c9",X"21",X"00",X"00",X"c9",X"c9",X"41",X"44", -- 1e88
  X"43",X"00",X"41",X"44",X"44",X"00",X"43",X"43", -- 1e90
  X"00",X"44",X"41",X"41",X"00",X"44",X"41",X"44", -- 1e98
  X"00",X"21",X"04",X"00",X"39",X"54",X"5d",X"cd", -- 1ea0
  X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"e5", -- 1ea8
  X"21",X"04",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 1eb0
  X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"cd",X"40", -- 1eb8
  X"2f",X"d1",X"7d",X"12",X"7c",X"b5",X"ca",X"cc", -- 1ec0
  X"1e",X"c3",X"a1",X"1e",X"c9",X"21",X"04",X"00", -- 1ec8
  X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"eb", -- 1ed0
  X"c1",X"e1",X"e5",X"c5",X"cd",X"40",X"2f",X"cd", -- 1ed8
  X"a8",X"2f",X"7c",X"b5",X"ca",X"17",X"1f",X"21", -- 1ee0
  X"04",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40", -- 1ee8
  X"2f",X"7c",X"b5",X"c2",X"fa",X"1e",X"21",X"00", -- 1ef0
  X"00",X"c9",X"21",X"04",X"00",X"39",X"54",X"5d", -- 1ef8
  X"cd",X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"21", -- 1f00
  X"02",X"00",X"39",X"54",X"5d",X"cd",X"4d",X"2f", -- 1f08
  X"23",X"cd",X"8d",X"2f",X"c3",X"cd",X"1e",X"21", -- 1f10
  X"04",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40", -- 1f18
  X"2f",X"eb",X"c1",X"e1",X"e5",X"c5",X"cd",X"40", -- 1f20
  X"2f",X"cd",X"04",X"30",X"c9",X"21",X"f3",X"ff", -- 1f28
  X"39",X"f9",X"21",X"0b",X"00",X"39",X"eb",X"21", -- 1f30
  X"00",X"00",X"cd",X"8d",X"2f",X"21",X"0b",X"00", -- 1f38
  X"39",X"cd",X"4d",X"2f",X"eb",X"21",X"08",X"00", -- 1f40
  X"cd",X"c8",X"2f",X"7c",X"b5",X"ca",X"7a",X"1f", -- 1f48
  X"c3",X"64",X"1f",X"21",X"0b",X"00",X"39",X"54", -- 1f50
  X"5d",X"cd",X"4d",X"2f",X"23",X"cd",X"8d",X"2f", -- 1f58
  X"2b",X"c3",X"3d",X"1f",X"21",X"00",X"00",X"39", -- 1f60
  X"eb",X"21",X"0b",X"00",X"39",X"cd",X"4d",X"2f", -- 1f68
  X"19",X"eb",X"21",X"20",X"00",X"7d",X"12",X"c3", -- 1f70
  X"53",X"1f",X"21",X"08",X"00",X"39",X"e5",X"21", -- 1f78
  X"13",X"00",X"39",X"cd",X"4d",X"2f",X"eb",X"21", -- 1f80
  X"00",X"00",X"cd",X"c2",X"2f",X"7c",X"b5",X"ca", -- 1f88
  X"98",X"1f",X"21",X"2b",X"00",X"c3",X"9b",X"1f", -- 1f90
  X"21",X"2d",X"00",X"d1",X"7d",X"12",X"21",X"0b", -- 1f98
  X"00",X"39",X"eb",X"21",X"07",X"00",X"cd",X"8d", -- 1fa0
  X"2f",X"21",X"00",X"00",X"39",X"eb",X"21",X"0b", -- 1fa8
  X"00",X"39",X"cd",X"4d",X"2f",X"19",X"e5",X"21", -- 1fb0
  X"13",X"00",X"39",X"cd",X"4d",X"2f",X"eb",X"21", -- 1fb8
  X"0a",X"00",X"cd",X"ab",X"2e",X"eb",X"11",X"30", -- 1fc0
  X"00",X"19",X"d1",X"7d",X"12",X"21",X"11",X"00", -- 1fc8
  X"39",X"e5",X"21",X"13",X"00",X"39",X"cd",X"4d", -- 1fd0
  X"2f",X"eb",X"21",X"0a",X"00",X"cd",X"ab",X"2e", -- 1fd8
  X"d1",X"cd",X"8d",X"2f",X"21",X"0b",X"00",X"39", -- 1fe0
  X"54",X"5d",X"cd",X"4d",X"2f",X"2b",X"cd",X"8d", -- 1fe8
  X"2f",X"23",X"21",X"11",X"00",X"39",X"cd",X"4d", -- 1ff0
  X"2f",X"af",X"b4",X"fa",X"05",X"20",X"b5",X"ca", -- 1ff8
  X"05",X"20",X"c3",X"a9",X"1f",X"21",X"00",X"00", -- 2000
  X"39",X"eb",X"21",X"0b",X"00",X"39",X"cd",X"4d", -- 2008
  X"2f",X"19",X"eb",X"21",X"08",X"00",X"39",X"cd", -- 2010
  X"40",X"2f",X"7d",X"12",X"21",X"09",X"00",X"39", -- 2018
  X"eb",X"21",X"00",X"00",X"cd",X"8d",X"2f",X"21", -- 2020
  X"0b",X"00",X"39",X"cd",X"4d",X"2f",X"eb",X"21", -- 2028
  X"08",X"00",X"cd",X"c8",X"2f",X"7c",X"b5",X"ca", -- 2030
  X"71",X"20",X"21",X"0f",X"00",X"39",X"cd",X"4d", -- 2038
  X"2f",X"e5",X"21",X"0b",X"00",X"39",X"54",X"5d", -- 2040
  X"cd",X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b", -- 2048
  X"d1",X"19",X"e5",X"21",X"02",X"00",X"39",X"e5", -- 2050
  X"21",X"0f",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 2058
  X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"d1",X"19", -- 2060
  X"cd",X"40",X"2f",X"d1",X"7d",X"12",X"c3",X"27", -- 2068
  X"20",X"21",X"0f",X"00",X"39",X"cd",X"4d",X"2f", -- 2070
  X"eb",X"21",X"09",X"00",X"39",X"cd",X"4d",X"2f", -- 2078
  X"19",X"eb",X"21",X"00",X"00",X"7d",X"12",X"21", -- 2080
  X"0d",X"00",X"39",X"f9",X"c9",X"c5",X"c5",X"21", -- 2088
  X"00",X"00",X"39",X"e5",X"21",X"04",X"00",X"39", -- 2090
  X"eb",X"21",X"00",X"00",X"cd",X"8d",X"2f",X"d1", -- 2098
  X"cd",X"8d",X"2f",X"21",X"06",X"00",X"39",X"cd", -- 20a0
  X"4d",X"2f",X"cd",X"40",X"2f",X"eb",X"21",X"2b", -- 20a8
  X"00",X"cd",X"a8",X"2f",X"7c",X"b5",X"c2",X"d5", -- 20b0
  X"20",X"21",X"06",X"00",X"39",X"cd",X"4d",X"2f", -- 20b8
  X"cd",X"40",X"2f",X"eb",X"21",X"2d",X"00",X"cd", -- 20c0
  X"a8",X"2f",X"7c",X"b5",X"c2",X"d5",X"20",X"21", -- 20c8
  X"00",X"00",X"c3",X"d8",X"20",X"21",X"01",X"00", -- 20d0
  X"7c",X"b5",X"ca",X"07",X"21",X"21",X"06",X"00", -- 20d8
  X"39",X"54",X"5d",X"cd",X"4d",X"2f",X"23",X"cd", -- 20e0
  X"8d",X"2f",X"2b",X"cd",X"40",X"2f",X"eb",X"21", -- 20e8
  X"2d",X"00",X"cd",X"a8",X"2f",X"7c",X"b5",X"ca", -- 20f0
  X"07",X"21",X"21",X"00",X"00",X"39",X"eb",X"e1", -- 20f8
  X"e5",X"cd",X"0b",X"30",X"cd",X"8d",X"2f",X"21", -- 2100
  X"06",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40", -- 2108
  X"2f",X"7c",X"b5",X"ca",X"4a",X"21",X"21",X"02", -- 2110
  X"00",X"39",X"e5",X"21",X"04",X"00",X"39",X"cd", -- 2118
  X"4d",X"2f",X"11",X"0a",X"00",X"cd",X"8b",X"2e", -- 2120
  X"e5",X"21",X"0a",X"00",X"39",X"54",X"5d",X"cd", -- 2128
  X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"cd", -- 2130
  X"40",X"2f",X"d1",X"19",X"eb",X"21",X"30",X"00", -- 2138
  X"cd",X"04",X"30",X"d1",X"cd",X"8d",X"2f",X"c3", -- 2140
  X"07",X"21",X"e1",X"e5",X"7c",X"b5",X"ca",X"5b", -- 2148
  X"21",X"c1",X"e1",X"e5",X"c5",X"cd",X"0b",X"30", -- 2150
  X"c1",X"c1",X"c9",X"c1",X"e1",X"e5",X"c5",X"c1", -- 2158
  X"c1",X"c9",X"c5",X"21",X"01",X"00",X"39",X"eb", -- 2160
  X"21",X"00",X"00",X"7d",X"12",X"21",X"04",X"00", -- 2168
  X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"7c", -- 2170
  X"b5",X"ca",X"92",X"22",X"21",X"04",X"00",X"39", -- 2178
  X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"eb",X"21", -- 2180
  X"30",X"00",X"cd",X"c2",X"2f",X"7c",X"b5",X"ca", -- 2188
  X"ae",X"21",X"21",X"04",X"00",X"39",X"cd",X"4d", -- 2190
  X"2f",X"cd",X"40",X"2f",X"eb",X"21",X"39",X"00", -- 2198
  X"cd",X"bb",X"2f",X"7c",X"b5",X"ca",X"ae",X"21", -- 21a0
  X"21",X"01",X"00",X"c3",X"b1",X"21",X"21",X"00", -- 21a8
  X"00",X"7c",X"b5",X"ca",X"c3",X"21",X"21",X"00", -- 21b0
  X"00",X"39",X"eb",X"21",X"30",X"00",X"7d",X"12", -- 21b8
  X"c3",X"54",X"22",X"21",X"04",X"00",X"39",X"cd", -- 21c0
  X"4d",X"2f",X"cd",X"40",X"2f",X"eb",X"21",X"41", -- 21c8
  X"00",X"cd",X"c2",X"2f",X"7c",X"b5",X"ca",X"f5", -- 21d0
  X"21",X"21",X"04",X"00",X"39",X"cd",X"4d",X"2f", -- 21d8
  X"cd",X"40",X"2f",X"eb",X"21",X"46",X"00",X"cd", -- 21e0
  X"bb",X"2f",X"7c",X"b5",X"ca",X"f5",X"21",X"21", -- 21e8
  X"01",X"00",X"c3",X"f8",X"21",X"21",X"00",X"00", -- 21f0
  X"7c",X"b5",X"ca",X"0a",X"22",X"21",X"00",X"00", -- 21f8
  X"39",X"eb",X"21",X"37",X"00",X"7d",X"12",X"c3", -- 2200
  X"54",X"22",X"21",X"04",X"00",X"39",X"cd",X"4d", -- 2208
  X"2f",X"cd",X"40",X"2f",X"eb",X"21",X"61",X"00", -- 2210
  X"cd",X"c2",X"2f",X"7c",X"b5",X"ca",X"3c",X"22", -- 2218
  X"21",X"04",X"00",X"39",X"cd",X"4d",X"2f",X"cd", -- 2220
  X"40",X"2f",X"eb",X"21",X"66",X"00",X"cd",X"bb", -- 2228
  X"2f",X"7c",X"b5",X"ca",X"3c",X"22",X"21",X"01", -- 2230
  X"00",X"c3",X"3f",X"22",X"21",X"00",X"00",X"7c", -- 2238
  X"b5",X"ca",X"51",X"22",X"21",X"00",X"00",X"39", -- 2240
  X"eb",X"21",X"57",X"00",X"7d",X"12",X"c3",X"54", -- 2248
  X"22",X"c3",X"92",X"22",X"21",X"01",X"00",X"39", -- 2250
  X"e5",X"21",X"03",X"00",X"39",X"cd",X"40",X"2f", -- 2258
  X"eb",X"21",X"04",X"00",X"cd",X"31",X"2f",X"eb", -- 2260
  X"21",X"06",X"00",X"39",X"cd",X"4d",X"2f",X"cd", -- 2268
  X"40",X"2f",X"19",X"eb",X"21",X"02",X"00",X"39", -- 2270
  X"cd",X"40",X"2f",X"cd",X"04",X"30",X"d1",X"7d", -- 2278
  X"12",X"21",X"04",X"00",X"39",X"54",X"5d",X"cd", -- 2280
  X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"c3", -- 2288
  X"6d",X"21",X"21",X"01",X"00",X"39",X"cd",X"40", -- 2290
  X"2f",X"c1",X"c9",X"c5",X"c5",X"21",X"02",X"00", -- 2298
  X"39",X"eb",X"21",X"00",X"00",X"cd",X"8d",X"2f", -- 22a0
  X"21",X"06",X"00",X"39",X"cd",X"4d",X"2f",X"cd", -- 22a8
  X"40",X"2f",X"7c",X"b5",X"ca",X"ce",X"23",X"21", -- 22b0
  X"06",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40", -- 22b8
  X"2f",X"eb",X"21",X"30",X"00",X"cd",X"c2",X"2f", -- 22c0
  X"7c",X"b5",X"ca",X"e9",X"22",X"21",X"06",X"00", -- 22c8
  X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"eb", -- 22d0
  X"21",X"39",X"00",X"cd",X"bb",X"2f",X"7c",X"b5", -- 22d8
  X"ca",X"e9",X"22",X"21",X"01",X"00",X"c3",X"ec", -- 22e0
  X"22",X"21",X"00",X"00",X"7c",X"b5",X"ca",X"ff", -- 22e8
  X"22",X"21",X"00",X"00",X"39",X"eb",X"21",X"30", -- 22f0
  X"00",X"cd",X"8d",X"2f",X"c3",X"92",X"23",X"21", -- 22f8
  X"06",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40", -- 2300
  X"2f",X"eb",X"21",X"41",X"00",X"cd",X"c2",X"2f", -- 2308
  X"7c",X"b5",X"ca",X"31",X"23",X"21",X"06",X"00", -- 2310
  X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"eb", -- 2318
  X"21",X"46",X"00",X"cd",X"bb",X"2f",X"7c",X"b5", -- 2320
  X"ca",X"31",X"23",X"21",X"01",X"00",X"c3",X"34", -- 2328
  X"23",X"21",X"00",X"00",X"7c",X"b5",X"ca",X"47", -- 2330
  X"23",X"21",X"00",X"00",X"39",X"eb",X"21",X"37", -- 2338
  X"00",X"cd",X"8d",X"2f",X"c3",X"92",X"23",X"21", -- 2340
  X"06",X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40", -- 2348
  X"2f",X"eb",X"21",X"61",X"00",X"cd",X"c2",X"2f", -- 2350
  X"7c",X"b5",X"ca",X"79",X"23",X"21",X"06",X"00", -- 2358
  X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f",X"eb", -- 2360
  X"21",X"66",X"00",X"cd",X"bb",X"2f",X"7c",X"b5", -- 2368
  X"ca",X"79",X"23",X"21",X"01",X"00",X"c3",X"7c", -- 2370
  X"23",X"21",X"00",X"00",X"7c",X"b5",X"ca",X"8f", -- 2378
  X"23",X"21",X"00",X"00",X"39",X"eb",X"21",X"57", -- 2380
  X"00",X"cd",X"8d",X"2f",X"c3",X"92",X"23",X"c3", -- 2388
  X"ce",X"23",X"21",X"02",X"00",X"39",X"e5",X"21", -- 2390
  X"04",X"00",X"39",X"cd",X"4d",X"2f",X"eb",X"21", -- 2398
  X"04",X"00",X"cd",X"31",X"2f",X"eb",X"21",X"08", -- 23a0
  X"00",X"39",X"cd",X"4d",X"2f",X"cd",X"40",X"2f", -- 23a8
  X"19",X"eb",X"c1",X"e1",X"e5",X"c5",X"cd",X"04", -- 23b0
  X"30",X"d1",X"cd",X"8d",X"2f",X"21",X"06",X"00", -- 23b8
  X"39",X"54",X"5d",X"cd",X"4d",X"2f",X"23",X"cd", -- 23c0
  X"8d",X"2f",X"2b",X"c3",X"a8",X"22",X"c1",X"e1", -- 23c8
  X"e5",X"c5",X"c1",X"c1",X"c9",X"21",X"e0",X"23", -- 23d0
  X"e5",X"3e",X"01",X"cd",X"68",X"25",X"c1",X"c9", -- 23d8
  X"0d",X"0a",X"00",X"21",X"f8",X"ff",X"39",X"f9", -- 23e0
  X"21",X"00",X"00",X"39",X"eb",X"21",X"03",X"00", -- 23e8
  X"cd",X"8d",X"2f",X"e1",X"e5",X"af",X"b4",X"fa", -- 23f0
  X"89",X"24",X"c3",X"0e",X"24",X"21",X"00",X"00", -- 23f8
  X"39",X"54",X"5d",X"cd",X"4d",X"2f",X"2b",X"cd", -- 2400
  X"8d",X"2f",X"23",X"c3",X"f3",X"23",X"21",X"07", -- 2408
  X"00",X"39",X"e5",X"21",X"0c",X"00",X"39",X"cd", -- 2410
  X"4d",X"2f",X"eb",X"21",X"0f",X"00",X"cd",X"a1", -- 2418
  X"2f",X"d1",X"7d",X"12",X"21",X"0a",X"00",X"39", -- 2420
  X"e5",X"21",X"0c",X"00",X"39",X"cd",X"4d",X"2f", -- 2428
  X"eb",X"21",X"04",X"00",X"cd",X"23",X"2f",X"eb", -- 2430
  X"21",X"ff",X"0f",X"cd",X"a1",X"2f",X"d1",X"cd", -- 2438
  X"8d",X"2f",X"21",X"07",X"00",X"39",X"cd",X"40", -- 2440
  X"2f",X"eb",X"21",X"0a",X"00",X"cd",X"c8",X"2f", -- 2448
  X"7c",X"b5",X"ca",X"6f",X"24",X"21",X"02",X"00", -- 2450
  X"39",X"eb",X"e1",X"e5",X"19",X"e5",X"21",X"09", -- 2458
  X"00",X"39",X"cd",X"40",X"2f",X"11",X"30",X"00", -- 2460
  X"19",X"d1",X"7d",X"12",X"c3",X"86",X"24",X"21", -- 2468
  X"02",X"00",X"39",X"eb",X"e1",X"e5",X"19",X"e5", -- 2470
  X"21",X"09",X"00",X"39",X"cd",X"40",X"2f",X"11", -- 2478
  X"37",X"00",X"19",X"d1",X"7d",X"12",X"c3",X"fd", -- 2480
  X"23",X"21",X"02",X"00",X"39",X"11",X"04",X"00", -- 2488
  X"19",X"eb",X"21",X"00",X"00",X"7d",X"12",X"21", -- 2490
  X"02",X"00",X"39",X"e5",X"3e",X"01",X"cd",X"68", -- 2498
  X"25",X"c1",X"21",X"08",X"00",X"39",X"f9",X"c9", -- 24a0
  X"c5",X"c5",X"c5",X"21",X"00",X"00",X"39",X"eb", -- 24a8
  X"21",X"01",X"00",X"cd",X"8d",X"2f",X"e1",X"e5", -- 24b0
  X"af",X"b4",X"fa",X"4b",X"25",X"c3",X"d1",X"24", -- 24b8
  X"21",X"00",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 24c0
  X"2f",X"2b",X"cd",X"8d",X"2f",X"23",X"c3",X"b6", -- 24c8
  X"24",X"21",X"05",X"00",X"39",X"e5",X"21",X"0a", -- 24d0
  X"00",X"39",X"cd",X"40",X"2f",X"eb",X"21",X"0f", -- 24d8
  X"00",X"cd",X"a1",X"2f",X"d1",X"7d",X"12",X"21", -- 24e0
  X"08",X"00",X"39",X"e5",X"21",X"0a",X"00",X"39", -- 24e8
  X"cd",X"40",X"2f",X"eb",X"21",X"04",X"00",X"cd", -- 24f0
  X"23",X"2f",X"eb",X"21",X"ff",X"0f",X"cd",X"a1", -- 24f8
  X"2f",X"d1",X"7d",X"12",X"21",X"05",X"00",X"39", -- 2500
  X"cd",X"40",X"2f",X"eb",X"21",X"0a",X"00",X"cd", -- 2508
  X"c8",X"2f",X"7c",X"b5",X"ca",X"31",X"25",X"21", -- 2510
  X"02",X"00",X"39",X"eb",X"e1",X"e5",X"19",X"e5", -- 2518
  X"21",X"07",X"00",X"39",X"cd",X"40",X"2f",X"11", -- 2520
  X"30",X"00",X"19",X"d1",X"7d",X"12",X"c3",X"48", -- 2528
  X"25",X"21",X"02",X"00",X"39",X"eb",X"e1",X"e5", -- 2530
  X"19",X"e5",X"21",X"07",X"00",X"39",X"cd",X"40", -- 2538
  X"2f",X"11",X"37",X"00",X"19",X"d1",X"7d",X"12", -- 2540
  X"c3",X"c0",X"24",X"21",X"02",X"00",X"39",X"11", -- 2548
  X"02",X"00",X"19",X"eb",X"21",X"00",X"00",X"7d", -- 2550
  X"12",X"21",X"02",X"00",X"39",X"e5",X"3e",X"01", -- 2558
  X"cd",X"68",X"25",X"c1",X"c1",X"c1",X"c1",X"c9", -- 2560
  X"c1",X"e1",X"e5",X"c5",X"cd",X"40",X"2f",X"7c", -- 2568
  X"b5",X"ca",X"8f",X"25",X"21",X"02",X"00",X"39", -- 2570
  X"54",X"5d",X"cd",X"4d",X"2f",X"23",X"cd",X"8d", -- 2578
  X"2f",X"2b",X"cd",X"40",X"2f",X"e5",X"3e",X"01", -- 2580
  X"cd",X"b7",X"26",X"c1",X"c3",X"68",X"25",X"c9", -- 2588
  X"3b",X"c5",X"21",X"00",X"00",X"39",X"eb",X"21", -- 2590
  X"00",X"00",X"cd",X"8d",X"2f",X"21",X"02",X"00", -- 2598
  X"39",X"e5",X"af",X"cd",X"c1",X"26",X"d1",X"7d", -- 25a0
  X"12",X"eb",X"21",X"0d",X"00",X"cd",X"ae",X"2f", -- 25a8
  X"7c",X"b5",X"ca",X"94",X"26",X"21",X"02",X"00", -- 25b0
  X"39",X"cd",X"40",X"2f",X"eb",X"21",X"09",X"00", -- 25b8
  X"cd",X"a8",X"2f",X"7c",X"b5",X"ca",X"d2",X"25", -- 25c0
  X"21",X"02",X"00",X"39",X"eb",X"21",X"20",X"00", -- 25c8
  X"7d",X"12",X"21",X"02",X"00",X"39",X"cd",X"40", -- 25d0
  X"2f",X"eb",X"21",X"08",X"00",X"cd",X"a8",X"2f", -- 25d8
  X"7c",X"b5",X"ca",X"f8",X"25",X"d1",X"d5",X"21", -- 25e0
  X"00",X"00",X"cd",X"b4",X"2f",X"7c",X"b5",X"ca", -- 25e8
  X"f8",X"25",X"21",X"01",X"00",X"c3",X"fb",X"25", -- 25f0
  X"21",X"00",X"00",X"7c",X"b5",X"ca",X"2f",X"26", -- 25f8
  X"21",X"00",X"00",X"39",X"54",X"5d",X"cd",X"4d", -- 2600
  X"2f",X"2b",X"cd",X"8d",X"2f",X"23",X"21",X"08", -- 2608
  X"00",X"e5",X"3e",X"01",X"cd",X"b7",X"26",X"c1", -- 2610
  X"21",X"20",X"00",X"e5",X"3e",X"01",X"cd",X"b7", -- 2618
  X"26",X"c1",X"21",X"08",X"00",X"e5",X"3e",X"01", -- 2620
  X"cd",X"b7",X"26",X"c1",X"c3",X"91",X"26",X"21", -- 2628
  X"02",X"00",X"39",X"cd",X"40",X"2f",X"e5",X"3e", -- 2630
  X"01",X"cd",X"38",X"1c",X"c1",X"7c",X"b5",X"ca", -- 2638
  X"59",X"26",X"d1",X"d5",X"21",X"05",X"00",X"39", -- 2640
  X"cd",X"4d",X"2f",X"cd",X"c8",X"2f",X"7c",X"b5", -- 2648
  X"ca",X"59",X"26",X"21",X"01",X"00",X"c3",X"5c", -- 2650
  X"26",X"21",X"00",X"00",X"7c",X"b5",X"ca",X"91", -- 2658
  X"26",X"21",X"07",X"00",X"39",X"cd",X"4d",X"2f", -- 2660
  X"e5",X"21",X"02",X"00",X"39",X"54",X"5d",X"cd", -- 2668
  X"4d",X"2f",X"23",X"cd",X"8d",X"2f",X"2b",X"d1", -- 2670
  X"19",X"eb",X"21",X"02",X"00",X"39",X"cd",X"40", -- 2678
  X"2f",X"7d",X"12",X"21",X"02",X"00",X"39",X"cd", -- 2680
  X"40",X"2f",X"e5",X"3e",X"01",X"cd",X"b7",X"26", -- 2688
  X"c1",X"c3",X"9d",X"25",X"21",X"07",X"00",X"39", -- 2690
  X"cd",X"4d",X"2f",X"eb",X"e1",X"e5",X"19",X"eb", -- 2698
  X"21",X"00",X"00",X"7d",X"12",X"af",X"cd",X"d5", -- 26a0
  X"23",X"33",X"c1",X"c9",X"c1",X"d1",X"d5",X"c5", -- 26a8
  X"21",X"b6",X"26",X"e5",X"eb",X"e9",X"c9",X"c1", -- 26b0
  X"d1",X"d5",X"c5",X"0e",X"02",X"cd",X"05",X"00", -- 26b8
  X"c9",X"0e",X"06",X"1e",X"ff",X"cd",X"05",X"00", -- 26c0
  X"fe",X"00",X"ca",X"c1",X"26",X"fe",X"61",X"da", -- 26c8
  X"d9",X"26",X"fe",X"7b",X"d2",X"d9",X"26",X"e6", -- 26d0
  X"df",X"26",X"00",X"6f",X"c9",X"e1",X"c3",X"21", -- 26d8
  X"01",X"c9",X"3f",X"00",X"41",X"43",X"49",X"00", -- 26e0
  X"41",X"44",X"43",X"00",X"41",X"44",X"44",X"00", -- 26e8
  X"41",X"44",X"49",X"00",X"41",X"4e",X"41",X"00", -- 26f0
  X"41",X"4e",X"49",X"00",X"43",X"41",X"4c",X"4c", -- 26f8
  X"00",X"43",X"43",X"00",X"43",X"4d",X"00",X"43", -- 2700
  X"4d",X"41",X"00",X"43",X"4d",X"43",X"00",X"43", -- 2708
  X"4d",X"50",X"00",X"43",X"4e",X"5a",X"00",X"43", -- 2710
  X"50",X"00",X"43",X"50",X"45",X"00",X"43",X"50", -- 2718
  X"49",X"00",X"43",X"50",X"4f",X"00",X"43",X"5a", -- 2720
  X"00",X"44",X"41",X"41",X"00",X"44",X"41",X"44", -- 2728
  X"00",X"44",X"43",X"52",X"00",X"44",X"43",X"58", -- 2730
  X"00",X"44",X"49",X"00",X"45",X"49",X"00",X"48", -- 2738
  X"4c",X"54",X"00",X"49",X"4e",X"00",X"49",X"4e", -- 2740
  X"52",X"00",X"49",X"4e",X"58",X"00",X"4a",X"43", -- 2748
  X"00",X"4a",X"4e",X"43",X"00",X"4a",X"4d",X"00", -- 2750
  X"4a",X"4d",X"50",X"00",X"4a",X"4e",X"5a",X"00", -- 2758
  X"4a",X"50",X"00",X"4a",X"50",X"45",X"00",X"4a", -- 2760
  X"50",X"4f",X"00",X"4a",X"5a",X"00",X"4c",X"44", -- 2768
  X"41",X"00",X"4c",X"44",X"41",X"58",X"00",X"4c", -- 2770
  X"48",X"4c",X"44",X"00",X"4c",X"58",X"49",X"00", -- 2778
  X"4d",X"4f",X"56",X"00",X"4d",X"56",X"49",X"00", -- 2780
  X"4e",X"4f",X"50",X"00",X"4f",X"52",X"41",X"00", -- 2788
  X"4f",X"52",X"49",X"00",X"4f",X"55",X"54",X"00", -- 2790
  X"50",X"43",X"48",X"4c",X"00",X"50",X"4f",X"50", -- 2798
  X"00",X"50",X"55",X"53",X"48",X"00",X"52",X"41", -- 27a0
  X"4c",X"00",X"52",X"41",X"52",X"00",X"52",X"43", -- 27a8
  X"00",X"52",X"45",X"54",X"00",X"52",X"4c",X"43", -- 27b0
  X"00",X"52",X"4d",X"00",X"52",X"4e",X"43",X"00", -- 27b8
  X"52",X"4e",X"5a",X"00",X"52",X"50",X"00",X"52", -- 27c0
  X"50",X"45",X"00",X"52",X"50",X"4f",X"00",X"52", -- 27c8
  X"52",X"43",X"00",X"52",X"53",X"54",X"30",X"00", -- 27d0
  X"52",X"53",X"54",X"31",X"00",X"52",X"53",X"54", -- 27d8
  X"32",X"00",X"52",X"53",X"54",X"33",X"00",X"52", -- 27e0
  X"53",X"54",X"34",X"00",X"52",X"53",X"54",X"35", -- 27e8
  X"00",X"52",X"53",X"54",X"36",X"00",X"52",X"53", -- 27f0
  X"54",X"37",X"00",X"52",X"5a",X"00",X"53",X"42", -- 27f8
  X"42",X"00",X"53",X"42",X"49",X"00",X"53",X"48", -- 2800
  X"4c",X"44",X"00",X"53",X"50",X"48",X"4c",X"00", -- 2808
  X"53",X"54",X"41",X"00",X"53",X"54",X"41",X"58", -- 2810
  X"00",X"53",X"54",X"43",X"00",X"53",X"55",X"42", -- 2818
  X"00",X"53",X"55",X"49",X"00",X"58",X"43",X"48", -- 2820
  X"47",X"00",X"58",X"52",X"41",X"00",X"58",X"52", -- 2828
  X"49",X"00",X"58",X"54",X"48",X"4c",X"00",X"43", -- 2830
  X"4e",X"43",X"00",X"88",X"27",X"7c",X"27",X"14", -- 2838
  X"28",X"4a",X"27",X"46",X"27",X"31",X"27",X"84", -- 2840
  X"27",X"b5",X"27",X"e2",X"26",X"2d",X"27",X"72", -- 2848
  X"27",X"35",X"27",X"46",X"27",X"31",X"27",X"84", -- 2850
  X"27",X"cf",X"27",X"e2",X"26",X"7c",X"27",X"14", -- 2858
  X"28",X"4a",X"27",X"46",X"27",X"31",X"27",X"84", -- 2860
  X"27",X"a6",X"27",X"e2",X"26",X"2d",X"27",X"72", -- 2868
  X"27",X"35",X"27",X"46",X"27",X"31",X"27",X"84", -- 2870
  X"27",X"aa",X"27",X"e2",X"26",X"7c",X"27",X"06", -- 2878
  X"28",X"4a",X"27",X"46",X"27",X"31",X"27",X"84", -- 2880
  X"27",X"29",X"27",X"e2",X"26",X"2d",X"27",X"77", -- 2888
  X"27",X"35",X"27",X"46",X"27",X"31",X"27",X"84", -- 2890
  X"27",X"07",X"27",X"e2",X"26",X"7c",X"27",X"10", -- 2898
  X"28",X"4a",X"27",X"46",X"27",X"31",X"27",X"84", -- 28a0
  X"27",X"19",X"28",X"e2",X"26",X"2d",X"27",X"6e", -- 28a8
  X"27",X"35",X"27",X"46",X"27",X"31",X"27",X"84", -- 28b0
  X"27",X"0b",X"27",X"80",X"27",X"80",X"27",X"80", -- 28b8
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 28c0
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 28c8
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 28d0
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 28d8
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 28e0
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 28e8
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 28f0
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 28f8
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 2900
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 2908
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 2910
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 2918
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"3f", -- 2920
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 2928
  X"27",X"80",X"27",X"80",X"27",X"80",X"27",X"80", -- 2930
  X"27",X"80",X"27",X"ec",X"26",X"ec",X"26",X"ec", -- 2938
  X"26",X"ec",X"26",X"ec",X"26",X"ec",X"26",X"ec", -- 2940
  X"26",X"ec",X"26",X"e8",X"26",X"e8",X"26",X"e8", -- 2948
  X"26",X"e8",X"26",X"e8",X"26",X"e8",X"26",X"e8", -- 2950
  X"26",X"e8",X"26",X"1d",X"28",X"1d",X"28",X"1d", -- 2958
  X"28",X"1d",X"28",X"1d",X"28",X"1d",X"28",X"1d", -- 2960
  X"28",X"1d",X"28",X"fe",X"27",X"fe",X"27",X"fe", -- 2968
  X"27",X"fe",X"27",X"fe",X"27",X"fe",X"27",X"fe", -- 2970
  X"27",X"fe",X"27",X"f4",X"26",X"f4",X"26",X"f4", -- 2978
  X"26",X"f4",X"26",X"f4",X"26",X"f4",X"26",X"f4", -- 2980
  X"26",X"f4",X"26",X"2a",X"28",X"2a",X"28",X"2a", -- 2988
  X"28",X"2a",X"28",X"2a",X"28",X"2a",X"28",X"2a", -- 2990
  X"28",X"2a",X"28",X"8c",X"27",X"8c",X"27",X"8c", -- 2998
  X"27",X"8c",X"27",X"8c",X"27",X"8c",X"27",X"8c", -- 29a0
  X"27",X"8c",X"27",X"0f",X"27",X"0f",X"27",X"0f", -- 29a8
  X"27",X"0f",X"27",X"0f",X"27",X"0f",X"27",X"0f", -- 29b0
  X"27",X"0f",X"27",X"c0",X"27",X"9d",X"27",X"5c", -- 29b8
  X"27",X"58",X"27",X"13",X"27",X"a1",X"27",X"f0", -- 29c0
  X"26",X"d3",X"27",X"fb",X"27",X"b1",X"27",X"6b", -- 29c8
  X"27",X"e2",X"26",X"26",X"27",X"fc",X"26",X"e4", -- 29d0
  X"26",X"d8",X"27",X"bc",X"27",X"9d",X"27",X"51", -- 29d8
  X"27",X"94",X"27",X"37",X"28",X"a1",X"27",X"21", -- 29e0
  X"28",X"dd",X"27",X"ae",X"27",X"e2",X"26",X"4e", -- 29e8
  X"27",X"43",X"27",X"01",X"27",X"e2",X"26",X"02", -- 29f0
  X"28",X"e2",X"27",X"cb",X"27",X"9d",X"27",X"67", -- 29f8
  X"27",X"32",X"28",X"22",X"27",X"a1",X"27",X"f8", -- 2a00
  X"26",X"e7",X"27",X"c7",X"27",X"98",X"27",X"63", -- 2a08
  X"27",X"25",X"28",X"1a",X"27",X"e2",X"26",X"2e", -- 2a10
  X"28",X"ec",X"27",X"c4",X"27",X"9d",X"27",X"60", -- 2a18
  X"27",X"39",X"27",X"17",X"27",X"a1",X"27",X"90", -- 2a20
  X"27",X"f1",X"27",X"b9",X"27",X"0b",X"28",X"55", -- 2a28
  X"27",X"3c",X"27",X"04",X"27",X"e2",X"26",X"1e", -- 2a30
  X"27",X"f6",X"27",X"00",X"00",X"01",X"00",X"02", -- 2a38
  X"00",X"42",X"00",X"43",X"00",X"44",X"00",X"45", -- 2a40
  X"00",X"48",X"00",X"4c",X"00",X"4d",X"00",X"41", -- 2a48
  X"00",X"50",X"53",X"57",X"00",X"53",X"50",X"00", -- 2a50
  X"3b",X"2a",X"41",X"2a",X"41",X"2a",X"41",X"2a", -- 2a58
  X"41",X"2a",X"41",X"2a",X"41",X"2a",X"3b",X"2a", -- 2a60
  X"3b",X"2a",X"41",X"2a",X"41",X"2a",X"41",X"2a", -- 2a68
  X"43",X"2a",X"43",X"2a",X"43",X"2a",X"3b",X"2a", -- 2a70
  X"3b",X"2a",X"45",X"2a",X"45",X"2a",X"45",X"2a", -- 2a78
  X"45",X"2a",X"45",X"2a",X"45",X"2a",X"3b",X"2a", -- 2a80
  X"3b",X"2a",X"45",X"2a",X"45",X"2a",X"45",X"2a", -- 2a88
  X"47",X"2a",X"47",X"2a",X"47",X"2a",X"3b",X"2a", -- 2a90
  X"3b",X"2a",X"49",X"2a",X"3f",X"2a",X"49",X"2a", -- 2a98
  X"49",X"2a",X"49",X"2a",X"49",X"2a",X"3b",X"2a", -- 2aa0
  X"3b",X"2a",X"49",X"2a",X"3f",X"2a",X"49",X"2a", -- 2aa8
  X"4b",X"2a",X"4b",X"2a",X"4b",X"2a",X"3b",X"2a", -- 2ab0
  X"3b",X"2a",X"55",X"2a",X"3f",X"2a",X"55",X"2a", -- 2ab8
  X"4d",X"2a",X"4d",X"2a",X"4d",X"2a",X"3b",X"2a", -- 2ac0
  X"3b",X"2a",X"55",X"2a",X"3f",X"2a",X"55",X"2a", -- 2ac8
  X"4f",X"2a",X"4f",X"2a",X"4f",X"2a",X"3b",X"2a", -- 2ad0
  X"41",X"2a",X"41",X"2a",X"41",X"2a",X"41",X"2a", -- 2ad8
  X"41",X"2a",X"41",X"2a",X"41",X"2a",X"41",X"2a", -- 2ae0
  X"43",X"2a",X"43",X"2a",X"43",X"2a",X"43",X"2a", -- 2ae8
  X"43",X"2a",X"43",X"2a",X"43",X"2a",X"43",X"2a", -- 2af0
  X"45",X"2a",X"45",X"2a",X"45",X"2a",X"45",X"2a", -- 2af8
  X"45",X"2a",X"45",X"2a",X"45",X"2a",X"45",X"2a", -- 2b00
  X"47",X"2a",X"47",X"2a",X"47",X"2a",X"47",X"2a", -- 2b08
  X"47",X"2a",X"47",X"2a",X"47",X"2a",X"47",X"2a", -- 2b10
  X"49",X"2a",X"49",X"2a",X"49",X"2a",X"49",X"2a", -- 2b18
  X"49",X"2a",X"49",X"2a",X"49",X"2a",X"49",X"2a", -- 2b20
  X"4b",X"2a",X"4b",X"2a",X"4b",X"2a",X"4b",X"2a", -- 2b28
  X"4b",X"2a",X"4b",X"2a",X"4b",X"2a",X"4b",X"2a", -- 2b30
  X"4d",X"2a",X"4d",X"2a",X"4d",X"2a",X"4d",X"2a", -- 2b38
  X"4d",X"2a",X"4d",X"2a",X"3b",X"2a",X"4d",X"2a", -- 2b40
  X"4f",X"2a",X"4f",X"2a",X"4f",X"2a",X"4f",X"2a", -- 2b48
  X"4f",X"2a",X"4f",X"2a",X"4f",X"2a",X"4f",X"2a", -- 2b50
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2b58
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2b60
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2b68
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2b70
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2b78
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2b80
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2b88
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2b90
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2b98
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2ba0
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2ba8
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2bb0
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2bb8
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2bc0
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2bc8
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2bd0
  X"3b",X"2a",X"41",X"2a",X"3f",X"2a",X"3f",X"2a", -- 2bd8
  X"3f",X"2a",X"41",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2be0
  X"3b",X"2a",X"3b",X"2a",X"3f",X"2a",X"3f",X"2a", -- 2be8
  X"3f",X"2a",X"3f",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2bf0
  X"3b",X"2a",X"45",X"2a",X"3f",X"2a",X"3d",X"2a", -- 2bf8
  X"3f",X"2a",X"45",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2c00
  X"3b",X"2a",X"3b",X"2a",X"3f",X"2a",X"3d",X"2a", -- 2c08
  X"3f",X"2a",X"3f",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2c10
  X"3b",X"2a",X"49",X"2a",X"3f",X"2a",X"3b",X"2a", -- 2c18
  X"3f",X"2a",X"49",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2c20
  X"3b",X"2a",X"3b",X"2a",X"3f",X"2a",X"3b",X"2a", -- 2c28
  X"3f",X"2a",X"3f",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2c30
  X"3b",X"2a",X"51",X"2a",X"3f",X"2a",X"3b",X"2a", -- 2c38
  X"3f",X"2a",X"51",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2c40
  X"3b",X"2a",X"3b",X"2a",X"3f",X"2a",X"3b",X"2a", -- 2c48
  X"3f",X"2a",X"3f",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2c50
  X"3b",X"2a",X"3f",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2c58
  X"3b",X"2a",X"3b",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2c60
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2c68
  X"3b",X"2a",X"3b",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2c70
  X"3b",X"2a",X"3f",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2c78
  X"3b",X"2a",X"3b",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2c80
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2c88
  X"3b",X"2a",X"3b",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2c90
  X"3b",X"2a",X"3f",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2c98
  X"3b",X"2a",X"3b",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2ca0
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2ca8
  X"3b",X"2a",X"3b",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2cb0
  X"3b",X"2a",X"3f",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2cb8
  X"3b",X"2a",X"3b",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2cc0
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2cc8
  X"3b",X"2a",X"3b",X"2a",X"3d",X"2a",X"3b",X"2a", -- 2cd0
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2cd8
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2ce0
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2ce8
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2cf0
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2cf8
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2d00
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2d08
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2d10
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2d18
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2d20
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2d28
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2d30
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2d38
  X"49",X"2a",X"4b",X"2a",X"3b",X"2a",X"4f",X"2a", -- 2d40
  X"41",X"2a",X"43",X"2a",X"45",X"2a",X"47",X"2a", -- 2d48
  X"49",X"2a",X"4b",X"2a",X"4d",X"2a",X"4f",X"2a", -- 2d50
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2d58
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2d60
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2d68
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2d70
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2d78
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2d80
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2d88
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2d90
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2d98
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2da0
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2da8
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2db0
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2db8
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2dc0
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2dc8
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2dd0
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2dd8
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2de0
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2de8
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2df0
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2df8
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2e00
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2e08
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2e10
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2e18
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2e20
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2e28
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2e30
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2e38
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2e40
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2e48
  X"3b",X"2a",X"3b",X"2a",X"3b",X"2a",X"3b",X"2a", -- 2e50
  X"d1",X"c1",X"c5",X"d5",X"11",X"3b",X"28",X"26", -- 2e58
  X"00",X"69",X"29",X"19",X"5e",X"23",X"56",X"eb", -- 2e60
  X"c9",X"d1",X"c1",X"c5",X"d5",X"11",X"58",X"2a", -- 2e68
  X"26",X"00",X"69",X"29",X"19",X"5e",X"23",X"56", -- 2e70
  X"eb",X"c9",X"d1",X"c1",X"c5",X"d5",X"11",X"58", -- 2e78
  X"2c",X"26",X"00",X"69",X"29",X"19",X"5e",X"23", -- 2e80
  X"56",X"eb",X"c9",X"44",X"4d",X"21",X"00",X"00", -- 2e88
  X"79",X"0f",X"d2",X"96",X"2e",X"19",X"af",X"78", -- 2e90
  X"1f",X"47",X"79",X"1f",X"4f",X"b0",X"c8",X"af", -- 2e98
  X"7b",X"17",X"5f",X"7a",X"17",X"57",X"b3",X"c8", -- 2ea0
  X"c3",X"90",X"2e",X"44",X"4d",X"7a",X"a8",X"f5", -- 2ea8
  X"7a",X"b7",X"fc",X"ec",X"2e",X"78",X"b7",X"fc", -- 2eb0
  X"f4",X"2e",X"3e",X"10",X"f5",X"eb",X"11",X"00", -- 2eb8
  X"00",X"29",X"cd",X"fc",X"2e",X"ca",X"d8",X"2e", -- 2ec0
  X"cd",X"04",X"2f",X"fa",X"d8",X"2e",X"7d",X"f6", -- 2ec8
  X"01",X"6f",X"7b",X"91",X"5f",X"7a",X"98",X"57", -- 2ed0
  X"f1",X"3d",X"ca",X"e1",X"2e",X"f5",X"c3",X"c1", -- 2ed8
  X"2e",X"f1",X"f0",X"cd",X"ec",X"2e",X"eb",X"cd", -- 2ee0
  X"ec",X"2e",X"eb",X"c9",X"7a",X"2f",X"57",X"7b", -- 2ee8
  X"2f",X"5f",X"13",X"c9",X"78",X"2f",X"47",X"79", -- 2ef0
  X"2f",X"4f",X"03",X"c9",X"7b",X"17",X"5f",X"7a", -- 2ef8
  X"17",X"57",X"b3",X"c9",X"7b",X"91",X"7a",X"98", -- 2f00
  X"c9",X"eb",X"e1",X"4e",X"23",X"46",X"23",X"78", -- 2f08
  X"b1",X"ca",X"22",X"2f",X"7e",X"23",X"bb",X"7e", -- 2f10
  X"23",X"c2",X"0b",X"2f",X"ba",X"c2",X"0b",X"2f", -- 2f18
  X"60",X"69",X"e9",X"eb",X"1d",X"f8",X"7c",X"17", -- 2f20
  X"7c",X"1f",X"67",X"7d",X"1f",X"6f",X"c3",X"24", -- 2f28
  X"2f",X"eb",X"1d",X"f8",X"29",X"c3",X"32",X"2f", -- 2f30
  X"e9",X"19",X"c3",X"40",X"2f",X"23",X"23",X"39", -- 2f38
  X"7e",X"6f",X"07",X"9f",X"67",X"c9",X"19",X"c3", -- 2f40
  X"4d",X"2f",X"23",X"23",X"39",X"7e",X"23",X"66", -- 2f48
  X"6f",X"c9",X"23",X"23",X"39",X"54",X"5d",X"cd", -- 2f50
  X"40",X"2f",X"2b",X"7d",X"12",X"c9",X"23",X"23", -- 2f58
  X"39",X"54",X"5d",X"cd",X"40",X"2f",X"23",X"7d", -- 2f60
  X"12",X"c9",X"19",X"c1",X"d1",X"c5",X"7d",X"12", -- 2f68
  X"c9",X"23",X"23",X"39",X"54",X"5d",X"cd",X"4d", -- 2f70
  X"2f",X"2b",X"c3",X"8d",X"2f",X"23",X"23",X"39", -- 2f78
  X"54",X"5d",X"cd",X"4d",X"2f",X"23",X"c3",X"8d", -- 2f80
  X"2f",X"19",X"c1",X"d1",X"c5",X"7d",X"12",X"13", -- 2f88
  X"7c",X"12",X"c9",X"7d",X"b3",X"6f",X"7c",X"b2", -- 2f90
  X"67",X"c9",X"7d",X"ab",X"6f",X"7c",X"aa",X"67", -- 2f98
  X"c9",X"7d",X"a3",X"6f",X"7c",X"a2",X"67",X"c9", -- 2fa0
  X"cd",X"ce",X"2f",X"c8",X"2b",X"c9",X"cd",X"ce", -- 2fa8
  X"2f",X"c0",X"2b",X"c9",X"eb",X"cd",X"ce",X"2f", -- 2fb0
  X"d8",X"2b",X"c9",X"cd",X"ce",X"2f",X"c8",X"d8", -- 2fb8
  X"2b",X"c9",X"cd",X"ce",X"2f",X"d0",X"2b",X"c9", -- 2fc0
  X"cd",X"ce",X"2f",X"d8",X"2b",X"c9",X"7c",X"ee", -- 2fc8
  X"80",X"67",X"7a",X"ee",X"80",X"bc",X"c2",X"db", -- 2fd0
  X"2f",X"7b",X"bd",X"21",X"01",X"00",X"c9",X"cd", -- 2fd8
  X"f9",X"2f",X"d0",X"2b",X"c9",X"cd",X"f9",X"2f", -- 2fe0
  X"d8",X"2b",X"c9",X"eb",X"cd",X"f9",X"2f",X"d8", -- 2fe8
  X"2b",X"c9",X"cd",X"f9",X"2f",X"c8",X"d8",X"2b", -- 2ff0
  X"c9",X"7a",X"bc",X"c2",X"00",X"30",X"7b",X"bd", -- 2ff8
  X"21",X"01",X"00",X"c9",X"7b",X"95",X"6f",X"7a", -- 3000
  X"9c",X"67",X"c9",X"cd",X"10",X"30",X"23",X"c9", -- 3008
  X"7c",X"2f",X"67",X"7d",X"2f",X"6f",X"c9",X"7c", -- 3010
  X"b5",X"c2",X"1f",X"30",X"2e",X"01",X"c9",X"21", -- 3018
  X"00",X"00",X"c9",X"00",X"00",X"00",X"00",X"00", -- 3020
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3028
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3030
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3038
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3040
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3048
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3050
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3058
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3060
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3068
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3070
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3078
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3080
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3088
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3090
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3098
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3100
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3108
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3110
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3118
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3120
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3128
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3130
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3138
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3140
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3148
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3150
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3158
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3160
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3168
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3170
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3178
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3180
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3188
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3190
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3198
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3200
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3208
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3210
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3218
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3220
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3228
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3230
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3238
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3240
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3248
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3250
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3258
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3260
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3268
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3270
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3278
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3280
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3288
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3290
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3298
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3300
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3308
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3310
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3318
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3320
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3328
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3330
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3338
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3340
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3348
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3350
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3358
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3360
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3368
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3370
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3378
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3380
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3388
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3390
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3398
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3400
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3408
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3410
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3418
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3420
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3428
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3430
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3438
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3440
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3448
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3450
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3458
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3460
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3468
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3470
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3478
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3480
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3488
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3490
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3498
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3500
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3508
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3510
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3518
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3520
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3528
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3530
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3538
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3540
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3548
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3550
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3558
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3560
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3568
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3570
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3578
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3580
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3588
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3590
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3598
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3600
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3608
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3610
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3618
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3620
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3628
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3630
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3638
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3640
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3648
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3650
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3658
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3660
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3668
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3670
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3678
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3680
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3688
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3690
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3698
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3700
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3708
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3710
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3718
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3720
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3728
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3730
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3738
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3740
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3748
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3750
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3758
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3760
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3768
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3770
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3778
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3780
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3788
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3790
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3798
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3800
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3808
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3810
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3818
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3820
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3828
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3830
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3838
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3840
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3848
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3850
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3858
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3860
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3868
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3870
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3878
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3880
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3888
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3890
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3898
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3900
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3908
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3910
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3918
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3920
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3928
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3930
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3938
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3940
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3948
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3950
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3958
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3960
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3968
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3970
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3978
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3980
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3988
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3990
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3998
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3aa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3aa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ab0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ab8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ac0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ac8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ad0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ad8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ae0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ae8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3af0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3af8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ba0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ba8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3be0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3be8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ca0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ca8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ce0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ce8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3da0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3da8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3db0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3db8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3de0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3de8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3df0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3df8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ea0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ea8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3eb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3eb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ec0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ec8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ed0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ed8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ee0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ee8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ef0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ef8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fe0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fe8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ff0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"  -- 3ff8
  );

end package obj_code_pkg;
