-------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
-------------------------------------------------------------------------------
-- Generated from "MSBAS80.BIN"
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Package with utility functions for handling SoC object code.
use work.mcu80_pkg.all;

package obj_code_pkg is

-- Object code initialization constant.
constant object_code : obj_code_t(0 to 16383) := (
  X"f3",X"c3",X"b9",X"00",X"00",X"00",X"00",X"00", -- 0000
  X"c3",X"a7",X"00",X"00",X"00",X"00",X"00",X"00", -- 0008
  X"c3",X"79",X"00",X"00",X"00",X"00",X"00",X"00", -- 0010
  X"c3",X"b3",X"00",X"00",X"00",X"00",X"00",X"00", -- 0018
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0020
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0028
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0030
  X"c3",X"3b",X"00",X"f5",X"e5",X"db",X"01",X"e6", -- 0038
  X"02",X"ca",X"75",X"00",X"db",X"00",X"f5",X"3a", -- 0040
  X"43",X"80",X"fe",X"3f",X"c2",X"53",X"00",X"f1", -- 0048
  X"c3",X"75",X"00",X"2a",X"3f",X"80",X"23",X"7d", -- 0050
  X"fe",X"3f",X"c2",X"60",X"00",X"21",X"00",X"80", -- 0058
  X"22",X"3f",X"80",X"f1",X"77",X"3a",X"43",X"80", -- 0060
  X"3c",X"32",X"43",X"80",X"fe",X"30",X"da",X"75", -- 0068
  X"00",X"3e",X"17",X"d3",X"01",X"e1",X"f1",X"fb", -- 0070
  X"c9",X"3a",X"43",X"80",X"fe",X"00",X"ca",X"79", -- 0078
  X"00",X"e5",X"2a",X"41",X"80",X"23",X"7d",X"fe", -- 0080
  X"3f",X"c2",X"8f",X"00",X"21",X"00",X"80",X"f3", -- 0088
  X"22",X"41",X"80",X"3a",X"43",X"80",X"3d",X"32", -- 0090
  X"43",X"80",X"fe",X"05",X"d2",X"a3",X"00",X"3e", -- 0098
  X"37",X"d3",X"01",X"7e",X"fb",X"e1",X"c9",X"f5", -- 00a0
  X"db",X"01",X"e6",X"01",X"ca",X"a8",X"00",X"f1", -- 00a8
  X"d3",X"00",X"c9",X"3a",X"43",X"80",X"fe",X"00", -- 00b0
  X"c9",X"21",X"ed",X"80",X"f9",X"21",X"00",X"80", -- 00b8
  X"22",X"3f",X"80",X"22",X"41",X"80",X"af",X"32", -- 00c0
  X"43",X"80",X"d3",X"01",X"d3",X"01",X"d3",X"01", -- 00c8
  X"3e",X"40",X"d3",X"01",X"00",X"00",X"3e",X"4e", -- 00d0
  X"d3",X"01",X"00",X"00",X"3e",X"37",X"d3",X"01", -- 00d8
  X"fb",X"c3",X"e4",X"00",X"c3",X"ea",X"00",X"c3", -- 00e0
  X"5f",X"01",X"c3",X"f1",X"00",X"b0",X"09",X"27", -- 00e8
  X"11",X"21",X"45",X"80",X"f9",X"c3",X"59",X"1d", -- 00f0
  X"11",X"cf",X"03",X"06",X"63",X"21",X"45",X"80", -- 00f8
  X"1a",X"77",X"23",X"13",X"05",X"c2",X"00",X"01", -- 0100
  X"f9",X"cd",X"d0",X"05",X"cd",X"a6",X"0b",X"32", -- 0108
  X"ef",X"80",X"32",X"3e",X"81",X"21",X"a2",X"81", -- 0110
  X"23",X"7c",X"b5",X"ca",X"27",X"01",X"7e",X"47", -- 0118
  X"2f",X"77",X"be",X"70",X"ca",X"18",X"01",X"2b", -- 0120
  X"11",X"a1",X"81",X"cd",X"66",X"07",X"da",X"68", -- 0128
  X"01",X"11",X"ce",X"ff",X"22",X"f4",X"80",X"19", -- 0130
  X"22",X"9f",X"80",X"cd",X"ab",X"05",X"2a",X"9f", -- 0138
  X"80",X"11",X"ef",X"ff",X"19",X"11",X"3e",X"81", -- 0140
  X"7d",X"93",X"6f",X"7c",X"9a",X"67",X"e5",X"21", -- 0148
  X"80",X"01",X"cd",X"45",X"12",X"e1",X"cd",X"ea", -- 0150
  X"18",X"21",X"71",X"01",X"cd",X"45",X"12",X"31", -- 0158
  X"ab",X"80",X"cd",X"d0",X"05",X"c3",X"e9",X"04", -- 0160
  X"21",X"bd",X"01",X"cd",X"45",X"12",X"c3",X"6e", -- 0168
  X"01",X"20",X"42",X"79",X"74",X"65",X"73",X"20", -- 0170
  X"66",X"72",X"65",X"65",X"0d",X"0a",X"00",X"00", -- 0178
  X"49",X"4e",X"54",X"45",X"4c",X"38",X"30",X"38", -- 0180
  X"30",X"20",X"42",X"41",X"53",X"49",X"43",X"20", -- 0188
  X"56",X"65",X"72",X"20",X"34",X"2e",X"37",X"62", -- 0190
  X"0d",X"0a",X"43",X"6f",X"70",X"79",X"72",X"69", -- 0198
  X"67",X"68",X"74",X"20",X"28",X"43",X"29",X"20", -- 01a0
  X"31",X"39",X"37",X"38",X"20",X"62",X"79",X"20", -- 01a8
  X"4d",X"69",X"63",X"72",X"6f",X"73",X"6f",X"66", -- 01b0
  X"74",X"0d",X"0a",X"00",X"00",X"4d",X"65",X"6d", -- 01b8
  X"6f",X"72",X"79",X"20",X"73",X"69",X"7a",X"65", -- 01c0
  X"20",X"6e",X"6f",X"74",X"20",X"65",X"6e",X"6f", -- 01c8
  X"75",X"67",X"68",X"0d",X"0a",X"54",X"68",X"65", -- 01d0
  X"20",X"73",X"79",X"73",X"74",X"65",X"6d",X"20", -- 01d8
  X"69",X"73",X"20",X"73",X"74",X"6f",X"70",X"70", -- 01e0
  X"65",X"64",X"2e",X"0d",X"0a",X"00",X"00",X"5f", -- 01e8
  X"17",X"23",X"18",X"75",X"17",X"48",X"80",X"05", -- 01f0
  X"11",X"8c",X"14",X"33",X"11",X"e9",X"19",X"c8", -- 01f8
  X"1a",X"04",X"16",X"37",X"1a",X"3d",X"1b",X"43", -- 0200
  X"1b",X"a4",X"1b",X"b9",X"1b",X"e0",X"14",X"26", -- 0208
  X"1c",X"96",X"80",X"b7",X"13",X"cf",X"11",X"51", -- 0210
  X"14",X"c6",X"13",X"d7",X"13",X"48",X"1c",X"e5", -- 0218
  X"1c",X"e7",X"13",X"17",X"14",X"21",X"14",X"c5", -- 0220
  X"4e",X"44",X"c6",X"4f",X"52",X"ce",X"45",X"58", -- 0228
  X"54",X"c4",X"41",X"54",X"41",X"c9",X"4e",X"50", -- 0230
  X"55",X"54",X"c4",X"49",X"4d",X"d2",X"45",X"41", -- 0238
  X"44",X"cc",X"45",X"54",X"c7",X"4f",X"54",X"4f", -- 0240
  X"d2",X"55",X"4e",X"c9",X"46",X"d2",X"45",X"53", -- 0248
  X"54",X"4f",X"52",X"45",X"c7",X"4f",X"53",X"55", -- 0250
  X"42",X"d2",X"45",X"54",X"55",X"52",X"4e",X"d2", -- 0258
  X"45",X"4d",X"d3",X"54",X"4f",X"50",X"cf",X"55", -- 0260
  X"54",X"cf",X"4e",X"ce",X"55",X"4c",X"4c",X"d7", -- 0268
  X"41",X"49",X"54",X"c4",X"45",X"46",X"d0",X"4f", -- 0270
  X"4b",X"45",X"c4",X"4f",X"4b",X"45",X"d3",X"43", -- 0278
  X"52",X"45",X"45",X"4e",X"cc",X"49",X"4e",X"45", -- 0280
  X"53",X"c3",X"4c",X"53",X"d7",X"49",X"44",X"54", -- 0288
  X"48",X"cd",X"4f",X"4e",X"49",X"54",X"4f",X"52", -- 0290
  X"d3",X"45",X"54",X"d2",X"45",X"53",X"45",X"54", -- 0298
  X"d0",X"52",X"49",X"4e",X"54",X"c3",X"4f",X"4e", -- 02a0
  X"54",X"cc",X"49",X"53",X"54",X"c3",X"4c",X"45", -- 02a8
  X"41",X"52",X"c3",X"4c",X"4f",X"41",X"44",X"c3", -- 02b0
  X"53",X"41",X"56",X"45",X"ce",X"45",X"57",X"d4", -- 02b8
  X"41",X"42",X"28",X"d4",X"4f",X"c6",X"4e",X"d3", -- 02c0
  X"50",X"43",X"28",X"d4",X"48",X"45",X"4e",X"ce", -- 02c8
  X"4f",X"54",X"d3",X"54",X"45",X"50",X"ab",X"ad", -- 02d0
  X"aa",X"af",X"de",X"c1",X"4e",X"44",X"cf",X"52", -- 02d8
  X"be",X"bd",X"bc",X"d3",X"47",X"4e",X"c9",X"4e", -- 02e0
  X"54",X"c1",X"42",X"53",X"d5",X"53",X"52",X"c6", -- 02e8
  X"52",X"45",X"c9",X"4e",X"50",X"d0",X"4f",X"53", -- 02f0
  X"d3",X"51",X"52",X"d2",X"4e",X"44",X"cc",X"4f", -- 02f8
  X"47",X"c5",X"58",X"50",X"c3",X"4f",X"53",X"d3", -- 0300
  X"49",X"4e",X"d4",X"41",X"4e",X"c1",X"54",X"4e", -- 0308
  X"d0",X"45",X"45",X"4b",X"c4",X"45",X"45",X"4b", -- 0310
  X"d0",X"4f",X"49",X"4e",X"54",X"cc",X"45",X"4e", -- 0318
  X"d3",X"54",X"52",X"24",X"d6",X"41",X"4c",X"c1", -- 0320
  X"53",X"43",X"c3",X"48",X"52",X"24",X"c8",X"45", -- 0328
  X"58",X"24",X"c2",X"49",X"4e",X"24",X"cc",X"45", -- 0330
  X"46",X"54",X"24",X"d2",X"49",X"47",X"48",X"54", -- 0338
  X"24",X"cd",X"49",X"44",X"24",X"80",X"48",X"09", -- 0340
  X"41",X"08",X"20",X"0d",X"95",X"0a",X"27",X"0c", -- 0348
  X"5d",X"0f",X"56",X"0c",X"ac",X"0a",X"52",X"0a", -- 0350
  X"35",X"0a",X"24",X"0b",X"0a",X"09",X"41",X"0a", -- 0358
  X"70",X"0a",X"97",X"0a",X"46",X"09",X"98",X"14", -- 0360
  X"06",X"0b",X"87",X"09",X"9e",X"14",X"3b",X"11", -- 0368
  X"e7",X"14",X"31",X"1c",X"97",X"0a",X"15",X"1c", -- 0370
  X"08",X"1c",X"0d",X"1c",X"56",X"1d",X"99",X"80", -- 0378
  X"9c",X"80",X"48",X"0b",X"74",X"09",X"b2",X"07", -- 0380
  X"ef",X"09",X"97",X"0a",X"97",X"0a",X"aa",X"05", -- 0388
  X"79",X"d1",X"18",X"79",X"05",X"15",X"7c",X"43", -- 0390
  X"16",X"7c",X"a4",X"16",X"7f",X"f2",X"19",X"50", -- 0398
  X"b6",X"0e",X"46",X"b5",X"0e",X"4e",X"46",X"53", -- 03a0
  X"4e",X"52",X"47",X"4f",X"44",X"46",X"43",X"4f", -- 03a8
  X"56",X"4f",X"4d",X"55",X"4c",X"42",X"53",X"44", -- 03b0
  X"44",X"2f",X"30",X"49",X"44",X"54",X"4d",X"4f", -- 03b8
  X"53",X"4c",X"53",X"53",X"54",X"43",X"4e",X"55", -- 03c0
  X"46",X"4d",X"4f",X"48",X"58",X"42",X"4e",X"c3", -- 03c8
  X"5f",X"01",X"c3",X"c5",X"09",X"d3",X"00",X"c9", -- 03d0
  X"d6",X"00",X"6f",X"7c",X"de",X"00",X"67",X"78", -- 03d8
  X"de",X"00",X"47",X"3e",X"00",X"c9",X"00",X"00", -- 03e0
  X"00",X"35",X"4a",X"ca",X"99",X"39",X"1c",X"76", -- 03e8
  X"98",X"22",X"95",X"b3",X"98",X"0a",X"dd",X"47", -- 03f0
  X"98",X"53",X"d1",X"99",X"99",X"0a",X"1a",X"9f", -- 03f8
  X"98",X"65",X"bc",X"cd",X"98",X"d6",X"77",X"3e", -- 0400
  X"98",X"52",X"c7",X"4f",X"80",X"db",X"00",X"c9", -- 0408
  X"01",X"ff",X"1c",X"00",X"00",X"14",X"00",X"14", -- 0410
  X"00",X"00",X"00",X"00",X"00",X"c3",X"e3",X"06", -- 0418
  X"c3",X"00",X"00",X"c3",X"00",X"00",X"c3",X"00", -- 0420
  X"00",X"a2",X"81",X"fe",X"ff",X"3f",X"81",X"20", -- 0428
  X"45",X"72",X"72",X"6f",X"72",X"00",X"20",X"69", -- 0430
  X"6e",X"20",X"00",X"4f",X"6b",X"0d",X"0a",X"00", -- 0438
  X"00",X"42",X"72",X"65",X"61",X"6b",X"00",X"21", -- 0440
  X"04",X"00",X"39",X"7e",X"23",X"fe",X"81",X"c0", -- 0448
  X"4e",X"23",X"46",X"23",X"e5",X"69",X"60",X"7a", -- 0450
  X"b3",X"eb",X"ca",X"61",X"04",X"eb",X"cd",X"66", -- 0458
  X"07",X"01",X"0d",X"00",X"e1",X"c8",X"09",X"c3", -- 0460
  X"4b",X"04",X"cd",X"84",X"04",X"c5",X"e3",X"c1", -- 0468
  X"cd",X"66",X"07",X"7e",X"02",X"c8",X"0b",X"2b", -- 0470
  X"c3",X"70",X"04",X"e5",X"2a",X"1f",X"81",X"06", -- 0478
  X"00",X"09",X"09",X"3e",X"e5",X"3e",X"d0",X"95", -- 0480
  X"6f",X"3e",X"ff",X"9c",X"da",X"93",X"04",X"67", -- 0488
  X"39",X"e1",X"d8",X"1e",X"0c",X"c3",X"b2",X"04", -- 0490
  X"2a",X"0e",X"81",X"22",X"a1",X"80",X"1e",X"02", -- 0498
  X"01",X"1e",X"14",X"01",X"1e",X"00",X"01",X"1e", -- 04a0
  X"12",X"01",X"1e",X"22",X"01",X"1e",X"0a",X"01", -- 04a8
  X"1e",X"18",X"cd",X"d0",X"05",X"32",X"8a",X"80", -- 04b0
  X"cd",X"99",X"0b",X"21",X"a5",X"03",X"57",X"3e", -- 04b8
  X"3f",X"cd",X"77",X"07",X"19",X"7e",X"cd",X"77", -- 04c0
  X"07",X"cd",X"fa",X"08",X"cd",X"77",X"07",X"21", -- 04c8
  X"2f",X"04",X"cd",X"45",X"12",X"2a",X"a1",X"80", -- 04d0
  X"11",X"fe",X"ff",X"cd",X"66",X"07",X"ca",X"f1", -- 04d8
  X"00",X"7c",X"a5",X"3c",X"c4",X"e2",X"18",X"3e", -- 04e0
  X"c1",X"af",X"32",X"8a",X"80",X"cd",X"99",X"0b", -- 04e8
  X"21",X"3b",X"04",X"cd",X"45",X"12",X"21",X"ff", -- 04f0
  X"ff",X"22",X"a1",X"80",X"cd",X"e3",X"06",X"da", -- 04f8
  X"f6",X"04",X"cd",X"fa",X"08",X"3c",X"3d",X"ca", -- 0500
  X"f6",X"04",X"f5",X"cd",X"ca",X"09",X"d5",X"cd", -- 0508
  X"fa",X"05",X"47",X"d1",X"f1",X"d2",X"da",X"08", -- 0510
  X"d5",X"c5",X"af",X"32",X"11",X"81",X"cd",X"fa", -- 0518
  X"08",X"b7",X"f5",X"cd",X"8a",X"05",X"da",X"2f", -- 0520
  X"05",X"f1",X"f5",X"ca",X"6b",X"0a",X"b7",X"c5", -- 0528
  X"d2",X"46",X"05",X"eb",X"2a",X"1b",X"81",X"1a", -- 0530
  X"02",X"03",X"13",X"cd",X"66",X"07",X"c2",X"37", -- 0538
  X"05",X"60",X"69",X"22",X"1b",X"81",X"d1",X"f1", -- 0540
  X"ca",X"6d",X"05",X"2a",X"1b",X"81",X"e3",X"c1", -- 0548
  X"09",X"e5",X"cd",X"6a",X"04",X"e1",X"22",X"1b", -- 0550
  X"81",X"eb",X"74",X"d1",X"23",X"23",X"73",X"23", -- 0558
  X"72",X"23",X"11",X"a6",X"80",X"1a",X"77",X"23", -- 0560
  X"13",X"b7",X"c2",X"65",X"05",X"cd",X"b6",X"05", -- 0568
  X"23",X"eb",X"62",X"6b",X"7e",X"23",X"b6",X"ca", -- 0570
  X"f6",X"04",X"23",X"23",X"23",X"af",X"be",X"23", -- 0578
  X"c2",X"7e",X"05",X"eb",X"73",X"23",X"72",X"c3", -- 0580
  X"72",X"05",X"2a",X"a3",X"80",X"44",X"4d",X"7e", -- 0588
  X"23",X"b6",X"2b",X"c8",X"23",X"23",X"7e",X"23", -- 0590
  X"66",X"6f",X"cd",X"66",X"07",X"60",X"69",X"7e", -- 0598
  X"23",X"66",X"6f",X"3f",X"c8",X"3f",X"d0",X"c3", -- 05a0
  X"8d",X"05",X"c0",X"2a",X"a3",X"80",X"af",X"77", -- 05a8
  X"23",X"77",X"23",X"22",X"1b",X"81",X"2a",X"a3", -- 05b0
  X"80",X"2b",X"22",X"13",X"81",X"2a",X"f4",X"80", -- 05b8
  X"22",X"08",X"81",X"af",X"cd",X"0a",X"09",X"2a", -- 05c0
  X"1b",X"81",X"22",X"1d",X"81",X"22",X"1f",X"81", -- 05c8
  X"c1",X"2a",X"9f",X"80",X"f9",X"21",X"f8",X"80", -- 05d0
  X"22",X"f6",X"80",X"af",X"6f",X"67",X"22",X"19", -- 05d8
  X"81",X"32",X"10",X"81",X"22",X"23",X"81",X"e5", -- 05e0
  X"c5",X"2a",X"13",X"81",X"c9",X"3e",X"3f",X"cd", -- 05e8
  X"77",X"07",X"3e",X"20",X"cd",X"77",X"07",X"c3", -- 05f0
  X"93",X"80",X"af",X"32",X"f3",X"80",X"0e",X"05", -- 05f8
  X"11",X"a6",X"80",X"7e",X"fe",X"20",X"ca",X"82", -- 0600
  X"06",X"47",X"fe",X"22",X"ca",X"a2",X"06",X"b7", -- 0608
  X"ca",X"a9",X"06",X"3a",X"f3",X"80",X"b7",X"7e", -- 0610
  X"c2",X"82",X"06",X"fe",X"3f",X"3e",X"9e",X"ca", -- 0618
  X"82",X"06",X"7e",X"fe",X"30",X"da",X"2d",X"06", -- 0620
  X"fe",X"3c",X"da",X"82",X"06",X"d5",X"11",X"26", -- 0628
  X"02",X"c5",X"01",X"7e",X"06",X"c5",X"06",X"7f", -- 0630
  X"7e",X"fe",X"61",X"da",X"46",X"06",X"fe",X"7b", -- 0638
  X"d2",X"46",X"06",X"e6",X"5f",X"77",X"4e",X"eb", -- 0640
  X"23",X"b6",X"f2",X"48",X"06",X"04",X"7e",X"e6", -- 0648
  X"7f",X"c8",X"b9",X"c2",X"48",X"06",X"eb",X"e5", -- 0650
  X"13",X"1a",X"b7",X"fa",X"7a",X"06",X"4f",X"78", -- 0658
  X"fe",X"88",X"c2",X"69",X"06",X"cd",X"fa",X"08", -- 0660
  X"2b",X"23",X"7e",X"fe",X"61",X"da",X"72",X"06", -- 0668
  X"e6",X"5f",X"b9",X"ca",X"58",X"06",X"e1",X"c3", -- 0670
  X"46",X"06",X"48",X"f1",X"eb",X"c9",X"eb",X"79", -- 0678
  X"c1",X"d1",X"23",X"12",X"13",X"0c",X"d6",X"3a", -- 0680
  X"ca",X"90",X"06",X"fe",X"49",X"c2",X"93",X"06", -- 0688
  X"32",X"f3",X"80",X"d6",X"54",X"c2",X"03",X"06", -- 0690
  X"47",X"7e",X"b7",X"ca",X"a9",X"06",X"b8",X"ca", -- 0698
  X"82",X"06",X"23",X"12",X"0c",X"13",X"c3",X"99", -- 06a0
  X"06",X"21",X"a5",X"80",X"12",X"13",X"12",X"13", -- 06a8
  X"12",X"c9",X"3a",X"89",X"80",X"b7",X"3e",X"00", -- 06b0
  X"32",X"89",X"80",X"c2",X"c6",X"06",X"05",X"ca", -- 06b8
  X"e3",X"06",X"cd",X"77",X"07",X"3e",X"05",X"2b", -- 06c0
  X"ca",X"da",X"06",X"7e",X"cd",X"77",X"07",X"c3", -- 06c8
  X"ec",X"06",X"05",X"2b",X"cd",X"77",X"07",X"c2", -- 06d0
  X"ec",X"06",X"cd",X"77",X"07",X"cd",X"a6",X"0b", -- 06d8
  X"c3",X"e3",X"06",X"21",X"a6",X"80",X"06",X"01", -- 06e0
  X"af",X"32",X"89",X"80",X"cd",X"a1",X"07",X"4f", -- 06e8
  X"fe",X"7f",X"ca",X"b2",X"06",X"3a",X"89",X"80", -- 06f0
  X"b7",X"ca",X"05",X"07",X"3e",X"00",X"cd",X"77", -- 06f8
  X"07",X"af",X"32",X"89",X"80",X"79",X"fe",X"07", -- 0700
  X"ca",X"49",X"07",X"fe",X"03",X"cc",X"a6",X"0b", -- 0708
  X"37",X"c8",X"fe",X"0d",X"ca",X"a1",X"0b",X"fe", -- 0710
  X"15",X"ca",X"dd",X"06",X"fe",X"40",X"ca",X"da", -- 0718
  X"06",X"fe",X"5f",X"ca",X"d2",X"06",X"fe",X"08", -- 0720
  X"ca",X"d2",X"06",X"fe",X"12",X"c2",X"44",X"07", -- 0728
  X"c5",X"d5",X"e5",X"36",X"00",X"cd",X"68",X"1d", -- 0730
  X"21",X"a6",X"80",X"cd",X"45",X"12",X"e1",X"d1", -- 0738
  X"c1",X"c3",X"ec",X"06",X"fe",X"20",X"da",X"ec", -- 0740
  X"06",X"78",X"fe",X"49",X"3e",X"07",X"d2",X"5e", -- 0748
  X"07",X"79",X"71",X"32",X"11",X"81",X"23",X"04", -- 0750
  X"cd",X"77",X"07",X"c3",X"ec",X"06",X"cd",X"77", -- 0758
  X"07",X"3e",X"08",X"c3",X"58",X"07",X"7c",X"92", -- 0760
  X"c0",X"7d",X"93",X"c9",X"7e",X"e3",X"be",X"23", -- 0768
  X"e3",X"ca",X"fa",X"08",X"c3",X"9e",X"04",X"f5", -- 0770
  X"3a",X"8a",X"80",X"b7",X"c2",X"7a",X"12",X"f1", -- 0778
  X"c5",X"f5",X"fe",X"20",X"da",X"9b",X"07",X"3a", -- 0780
  X"87",X"80",X"47",X"3a",X"f0",X"80",X"04",X"ca", -- 0788
  X"97",X"07",X"05",X"b8",X"cc",X"a6",X"0b",X"3c", -- 0790
  X"32",X"f0",X"80",X"f1",X"c1",X"cd",X"53",X"1d", -- 0798
  X"c9",X"cd",X"06",X"1c",X"e6",X"7f",X"fe",X"0f", -- 07a0
  X"c0",X"3a",X"8a",X"80",X"2f",X"32",X"8a",X"80", -- 07a8
  X"af",X"c9",X"cd",X"ca",X"09",X"c0",X"c1",X"cd", -- 07b0
  X"8a",X"05",X"c5",X"cd",X"08",X"08",X"e1",X"4e", -- 07b8
  X"23",X"46",X"23",X"78",X"b1",X"ca",X"e9",X"04", -- 07c0
  X"cd",X"11",X"08",X"cd",X"25",X"09",X"c5",X"cd", -- 07c8
  X"a6",X"0b",X"5e",X"23",X"56",X"23",X"e5",X"eb", -- 07d0
  X"cd",X"ea",X"18",X"3e",X"20",X"e1",X"cd",X"77", -- 07d8
  X"07",X"7e",X"b7",X"23",X"ca",X"be",X"07",X"f2", -- 07e0
  X"de",X"07",X"d6",X"7f",X"4f",X"11",X"27",X"02", -- 07e8
  X"1a",X"13",X"b7",X"f2",X"f0",X"07",X"0d",X"c2", -- 07f0
  X"f0",X"07",X"e6",X"7f",X"cd",X"77",X"07",X"1a", -- 07f8
  X"13",X"b7",X"f2",X"fa",X"07",X"c3",X"e1",X"07", -- 0800
  X"e5",X"2a",X"8d",X"80",X"22",X"8b",X"80",X"e1", -- 0808
  X"c9",X"e5",X"d5",X"2a",X"8b",X"80",X"11",X"ff", -- 0810
  X"ff",X"7b",X"8d",X"6f",X"7a",X"8c",X"67",X"22", -- 0818
  X"8b",X"80",X"d1",X"e1",X"f0",X"e5",X"2a",X"8d", -- 0820
  X"80",X"22",X"8b",X"80",X"cd",X"06",X"1c",X"fe", -- 0828
  X"03",X"ca",X"38",X"08",X"e1",X"c3",X"11",X"08", -- 0830
  X"2a",X"8d",X"80",X"22",X"8b",X"80",X"c3",X"62", -- 0838
  X"01",X"3e",X"64",X"32",X"10",X"81",X"cd",X"ac", -- 0840
  X"0a",X"c1",X"e5",X"cd",X"95",X"0a",X"22",X"0c", -- 0848
  X"81",X"21",X"02",X"00",X"39",X"cd",X"4b",X"04", -- 0850
  X"d1",X"c2",X"71",X"08",X"09",X"d5",X"2b",X"56", -- 0858
  X"2b",X"5e",X"23",X"23",X"e5",X"2a",X"0c",X"81", -- 0860
  X"cd",X"66",X"07",X"e1",X"c2",X"55",X"08",X"d1", -- 0868
  X"f9",X"eb",X"0e",X"08",X"cd",X"7b",X"04",X"e5", -- 0870
  X"2a",X"0c",X"81",X"e3",X"e5",X"2a",X"a1",X"80", -- 0878
  X"e3",X"cd",X"6e",X"0d",X"cd",X"6c",X"07",X"a6", -- 0880
  X"cd",X"6b",X"0d",X"e5",X"cd",X"9c",X"17",X"e1", -- 0888
  X"c5",X"d5",X"01",X"00",X"81",X"51",X"5a",X"7e", -- 0890
  X"fe",X"ab",X"3e",X"01",X"c2",X"ad",X"08",X"cd", -- 0898
  X"fa",X"08",X"cd",X"6b",X"0d",X"e5",X"cd",X"9c", -- 08a0
  X"17",X"cd",X"50",X"17",X"e1",X"c5",X"d5",X"f5", -- 08a8
  X"33",X"e5",X"2a",X"13",X"81",X"e3",X"06",X"81", -- 08b0
  X"c5",X"33",X"cd",X"25",X"09",X"22",X"13",X"81", -- 08b8
  X"7e",X"fe",X"3a",X"ca",X"da",X"08",X"b7",X"c2", -- 08c0
  X"9e",X"04",X"23",X"7e",X"23",X"b6",X"ca",X"50", -- 08c8
  X"09",X"23",X"5e",X"23",X"56",X"eb",X"22",X"a1", -- 08d0
  X"80",X"eb",X"cd",X"fa",X"08",X"11",X"ba",X"08", -- 08d8
  X"d5",X"c8",X"d6",X"80",X"da",X"ac",X"0a",X"fe", -- 08e0
  X"25",X"d2",X"9e",X"04",X"07",X"4f",X"06",X"00", -- 08e8
  X"eb",X"21",X"46",X"03",X"09",X"4e",X"23",X"46", -- 08f0
  X"c5",X"eb",X"23",X"7e",X"fe",X"3a",X"d0",X"fe", -- 08f8
  X"20",X"ca",X"fa",X"08",X"fe",X"30",X"3f",X"3c", -- 0900
  X"3d",X"c9",X"eb",X"2a",X"a3",X"80",X"ca",X"1f", -- 0908
  X"09",X"eb",X"cd",X"ca",X"09",X"e5",X"cd",X"8a", -- 0910
  X"05",X"60",X"69",X"d1",X"d2",X"6b",X"0a",X"2b", -- 0918
  X"22",X"21",X"81",X"eb",X"c9",X"df",X"c8",X"d7", -- 0920
  X"fe",X"1b",X"ca",X"41",X"09",X"fe",X"03",X"ca", -- 0928
  X"41",X"09",X"fe",X"13",X"c0",X"d7",X"fe",X"11", -- 0930
  X"c8",X"fe",X"03",X"ca",X"46",X"09",X"c3",X"35", -- 0938
  X"09",X"3e",X"ff",X"32",X"92",X"80",X"c0",X"f6", -- 0940
  X"c0",X"22",X"13",X"81",X"21",X"f6",X"ff",X"c1", -- 0948
  X"2a",X"a1",X"80",X"f5",X"7d",X"a4",X"3c",X"ca", -- 0950
  X"63",X"09",X"22",X"17",X"81",X"2a",X"13",X"81", -- 0958
  X"22",X"19",X"81",X"af",X"32",X"8a",X"80",X"cd", -- 0960
  X"99",X"0b",X"f1",X"21",X"41",X"04",X"c2",X"d2", -- 0968
  X"04",X"c3",X"e9",X"04",X"2a",X"19",X"81",X"7c", -- 0970
  X"b5",X"1e",X"20",X"ca",X"b2",X"04",X"eb",X"2a", -- 0978
  X"17",X"81",X"22",X"a1",X"80",X"eb",X"c9",X"cd", -- 0980
  X"cf",X"14",X"c0",X"32",X"86",X"80",X"c9",X"e5", -- 0988
  X"2a",X"8f",X"80",X"06",X"00",X"4f",X"09",X"22", -- 0990
  X"8f",X"80",X"e1",X"c9",X"7e",X"fe",X"41",X"d8", -- 0998
  X"fe",X"5b",X"3f",X"c9",X"cd",X"fa",X"08",X"cd", -- 09a0
  X"6b",X"0d",X"cd",X"50",X"17",X"fa",X"c5",X"09", -- 09a8
  X"3a",X"2c",X"81",X"fe",X"90",X"da",X"f8",X"17", -- 09b0
  X"01",X"80",X"90",X"11",X"00",X"00",X"e5",X"cd", -- 09b8
  X"cb",X"17",X"e1",X"51",X"c8",X"1e",X"08",X"c3", -- 09c0
  X"b2",X"04",X"2b",X"11",X"00",X"00",X"cd",X"fa", -- 09c8
  X"08",X"d0",X"e5",X"f5",X"21",X"98",X"19",X"cd", -- 09d0
  X"66",X"07",X"da",X"9e",X"04",X"62",X"6b",X"19", -- 09d8
  X"29",X"19",X"29",X"f1",X"d6",X"30",X"5f",X"16", -- 09e0
  X"00",X"19",X"eb",X"e1",X"c3",X"ce",X"09",X"ca", -- 09e8
  X"ba",X"05",X"cd",X"a7",X"09",X"2b",X"cd",X"fa", -- 09f0
  X"08",X"e5",X"2a",X"f4",X"80",X"ca",X"12",X"0a", -- 09f8
  X"e1",X"cd",X"6c",X"07",X"2c",X"d5",X"cd",X"a7", -- 0a00
  X"09",X"2b",X"cd",X"fa",X"08",X"c2",X"9e",X"04", -- 0a08
  X"e3",X"eb",X"7d",X"93",X"5f",X"7c",X"9a",X"57", -- 0a10
  X"da",X"93",X"04",X"e5",X"2a",X"1b",X"81",X"01", -- 0a18
  X"28",X"00",X"09",X"cd",X"66",X"07",X"d2",X"93", -- 0a20
  X"04",X"eb",X"22",X"9f",X"80",X"e1",X"22",X"f4", -- 0a28
  X"80",X"e1",X"c3",X"ba",X"05",X"ca",X"b6",X"05", -- 0a30
  X"cd",X"ba",X"05",X"01",X"ba",X"08",X"c3",X"51", -- 0a38
  X"0a",X"0e",X"03",X"cd",X"7b",X"04",X"c1",X"e5", -- 0a40
  X"e5",X"2a",X"a1",X"80",X"e3",X"3e",X"8c",X"f5", -- 0a48
  X"33",X"c5",X"cd",X"ca",X"09",X"cd",X"97",X"0a", -- 0a50
  X"e5",X"2a",X"a1",X"80",X"cd",X"66",X"07",X"e1", -- 0a58
  X"23",X"dc",X"8d",X"05",X"d4",X"8a",X"05",X"60", -- 0a60
  X"69",X"2b",X"d8",X"1e",X"0e",X"c3",X"b2",X"04", -- 0a68
  X"c0",X"16",X"ff",X"cd",X"47",X"04",X"f9",X"fe", -- 0a70
  X"8c",X"1e",X"04",X"c2",X"b2",X"04",X"e1",X"22", -- 0a78
  X"a1",X"80",X"23",X"7c",X"b5",X"c2",X"8f",X"0a", -- 0a80
  X"3a",X"11",X"81",X"b7",X"c2",X"e8",X"04",X"21", -- 0a88
  X"ba",X"08",X"e3",X"3e",X"e1",X"01",X"3a",X"0e", -- 0a90
  X"00",X"06",X"00",X"79",X"48",X"47",X"7e",X"b7", -- 0a98
  X"c8",X"b8",X"c8",X"23",X"fe",X"22",X"ca",X"9b", -- 0aa0
  X"0a",X"c3",X"9e",X"0a",X"cd",X"62",X"0f",X"cd", -- 0aa8
  X"6c",X"07",X"b4",X"d5",X"3a",X"f2",X"80",X"f5", -- 0ab0
  X"cd",X"7d",X"0d",X"f1",X"e3",X"22",X"13",X"81", -- 0ab8
  X"1f",X"cd",X"70",X"0d",X"ca",X"ff",X"0a",X"e5", -- 0ac0
  X"2a",X"29",X"81",X"e5",X"23",X"23",X"5e",X"23", -- 0ac8
  X"56",X"2a",X"a3",X"80",X"cd",X"66",X"07",X"d2", -- 0ad0
  X"ee",X"0a",X"2a",X"9f",X"80",X"cd",X"66",X"07", -- 0ad8
  X"d1",X"d2",X"f6",X"0a",X"21",X"04",X"81",X"cd", -- 0ae0
  X"66",X"07",X"d2",X"f6",X"0a",X"3e",X"d1",X"cd", -- 0ae8
  X"a6",X"13",X"eb",X"cd",X"df",X"11",X"cd",X"a6", -- 0af0
  X"13",X"e1",X"cd",X"ab",X"17",X"e1",X"c9",X"e5", -- 0af8
  X"cd",X"a8",X"17",X"d1",X"e1",X"c9",X"cd",X"cf", -- 0b00
  X"14",X"7e",X"47",X"fe",X"8c",X"ca",X"15",X"0b", -- 0b08
  X"cd",X"6c",X"07",X"88",X"2b",X"4b",X"0d",X"78", -- 0b10
  X"ca",X"e2",X"08",X"cd",X"cb",X"09",X"fe",X"2c", -- 0b18
  X"c0",X"c3",X"16",X"0b",X"cd",X"7d",X"0d",X"7e", -- 0b20
  X"fe",X"88",X"ca",X"32",X"0b",X"cd",X"6c",X"07", -- 0b28
  X"a9",X"2b",X"cd",X"6e",X"0d",X"cd",X"50",X"17", -- 0b30
  X"ca",X"97",X"0a",X"cd",X"fa",X"08",X"da",X"52", -- 0b38
  X"0a",X"c3",X"e1",X"08",X"2b",X"cd",X"fa",X"08", -- 0b40
  X"ca",X"a6",X"0b",X"c8",X"fe",X"a5",X"ca",X"d9", -- 0b48
  X"0b",X"fe",X"a8",X"ca",X"d9",X"0b",X"e5",X"fe", -- 0b50
  X"2c",X"ca",X"c2",X"0b",X"fe",X"3b",X"ca",X"fc", -- 0b58
  X"0b",X"c1",X"cd",X"7d",X"0d",X"e5",X"3a",X"f2", -- 0b60
  X"80",X"b7",X"c2",X"92",X"0b",X"cd",X"f5",X"18", -- 0b68
  X"cd",X"03",X"12",X"36",X"20",X"2a",X"29",X"81", -- 0b70
  X"34",X"2a",X"29",X"81",X"3a",X"87",X"80",X"47", -- 0b78
  X"04",X"ca",X"8e",X"0b",X"04",X"3a",X"f0",X"80", -- 0b80
  X"86",X"3d",X"b8",X"d4",X"a6",X"0b",X"cd",X"48", -- 0b88
  X"12",X"af",X"c4",X"48",X"12",X"e1",X"c3",X"44", -- 0b90
  X"0b",X"3a",X"f0",X"80",X"b7",X"c8",X"c3",X"a6", -- 0b98
  X"0b",X"36",X"00",X"21",X"a5",X"80",X"3e",X"0d", -- 0ba0
  X"cd",X"77",X"07",X"3e",X"0a",X"cd",X"77",X"07", -- 0ba8
  X"af",X"32",X"f0",X"80",X"3a",X"86",X"80",X"3d", -- 0bb0
  X"c8",X"f5",X"af",X"cd",X"77",X"07",X"f1",X"c3", -- 0bb8
  X"b7",X"0b",X"3a",X"88",X"80",X"47",X"3a",X"f0", -- 0bc0
  X"80",X"b8",X"d4",X"a6",X"0b",X"d2",X"fc",X"0b", -- 0bc8
  X"d6",X"0e",X"d2",X"d0",X"0b",X"2f",X"c3",X"f1", -- 0bd0
  X"0b",X"f5",X"cd",X"cc",X"14",X"cd",X"6c",X"07", -- 0bd8
  X"29",X"2b",X"f1",X"d6",X"a8",X"e5",X"ca",X"ec", -- 0be0
  X"0b",X"3a",X"f0",X"80",X"2f",X"83",X"d2",X"fc", -- 0be8
  X"0b",X"3c",X"47",X"3e",X"20",X"cd",X"77",X"07", -- 0bf0
  X"05",X"c2",X"f5",X"0b",X"e1",X"cd",X"fa",X"08", -- 0bf8
  X"c3",X"4b",X"0b",X"3f",X"52",X"65",X"64",X"6f", -- 0c00
  X"20",X"66",X"72",X"6f",X"6d",X"20",X"73",X"74", -- 0c08
  X"61",X"72",X"74",X"0d",X"0a",X"00",X"3a",X"12", -- 0c10
  X"81",X"b7",X"c2",X"98",X"04",X"c1",X"21",X"03", -- 0c18
  X"0c",X"cd",X"45",X"12",X"c3",X"e9",X"05",X"cd", -- 0c20
  X"b0",X"11",X"7e",X"fe",X"22",X"3e",X"00",X"32", -- 0c28
  X"8a",X"80",X"c2",X"41",X"0c",X"cd",X"04",X"12", -- 0c30
  X"cd",X"6c",X"07",X"3b",X"e5",X"cd",X"48",X"12", -- 0c38
  X"3e",X"e5",X"cd",X"ed",X"05",X"c1",X"da",X"4d", -- 0c40
  X"09",X"23",X"7e",X"b7",X"2b",X"c5",X"ca",X"94", -- 0c48
  X"0a",X"36",X"2c",X"c3",X"5b",X"0c",X"e5",X"2a", -- 0c50
  X"21",X"81",X"f6",X"af",X"32",X"12",X"81",X"e3", -- 0c58
  X"c3",X"67",X"0c",X"cd",X"6c",X"07",X"2c",X"cd", -- 0c60
  X"62",X"0f",X"e3",X"d5",X"7e",X"fe",X"2c",X"ca", -- 0c68
  X"8f",X"0c",X"3a",X"12",X"81",X"b7",X"c2",X"fc", -- 0c70
  X"0c",X"3e",X"3f",X"cd",X"77",X"07",X"cd",X"ed", -- 0c78
  X"05",X"d1",X"c1",X"da",X"4d",X"09",X"23",X"7e", -- 0c80
  X"b7",X"2b",X"c5",X"ca",X"94",X"0a",X"d5",X"3a", -- 0c88
  X"f2",X"80",X"b7",X"ca",X"b9",X"0c",X"cd",X"fa", -- 0c90
  X"08",X"57",X"47",X"fe",X"22",X"ca",X"ad",X"0c", -- 0c98
  X"3a",X"12",X"81",X"b7",X"57",X"ca",X"aa",X"0c", -- 0ca0
  X"16",X"3a",X"06",X"2c",X"2b",X"cd",X"07",X"12", -- 0ca8
  X"eb",X"21",X"c4",X"0c",X"e3",X"d5",X"c3",X"c7", -- 0cb0
  X"0a",X"cd",X"fa",X"08",X"cd",X"57",X"18",X"e3", -- 0cb8
  X"cd",X"a8",X"17",X"e1",X"2b",X"cd",X"fa",X"08", -- 0cc0
  X"ca",X"d0",X"0c",X"fe",X"2c",X"c2",X"16",X"0c", -- 0cc8
  X"e3",X"2b",X"cd",X"fa",X"08",X"c2",X"63",X"0c", -- 0cd0
  X"d1",X"3a",X"12",X"81",X"b7",X"eb",X"c2",X"20", -- 0cd8
  X"09",X"d5",X"b6",X"21",X"eb",X"0c",X"c4",X"45", -- 0ce0
  X"12",X"e1",X"c9",X"3f",X"45",X"78",X"74",X"72", -- 0ce8
  X"61",X"20",X"69",X"67",X"6e",X"6f",X"72",X"65", -- 0cf0
  X"64",X"0d",X"0a",X"00",X"cd",X"95",X"0a",X"b7", -- 0cf8
  X"c2",X"15",X"0d",X"23",X"7e",X"23",X"b6",X"1e", -- 0d00
  X"06",X"ca",X"b2",X"04",X"23",X"5e",X"23",X"56", -- 0d08
  X"eb",X"22",X"0e",X"81",X"eb",X"cd",X"fa",X"08", -- 0d10
  X"fe",X"83",X"c2",X"fc",X"0c",X"c3",X"8f",X"0c", -- 0d18
  X"11",X"00",X"00",X"c4",X"62",X"0f",X"22",X"13", -- 0d20
  X"81",X"cd",X"47",X"04",X"c2",X"a4",X"04",X"f9", -- 0d28
  X"d5",X"7e",X"23",X"f5",X"d5",X"cd",X"8e",X"17", -- 0d30
  X"e3",X"e5",X"cd",X"fb",X"14",X"e1",X"cd",X"a8", -- 0d38
  X"17",X"e1",X"cd",X"9f",X"17",X"e5",X"cd",X"cb", -- 0d40
  X"17",X"e1",X"c1",X"90",X"cd",X"9f",X"17",X"ca", -- 0d48
  X"5b",X"0d",X"eb",X"22",X"a1",X"80",X"69",X"60", -- 0d50
  X"c3",X"b6",X"08",X"f9",X"2a",X"13",X"81",X"7e", -- 0d58
  X"fe",X"2c",X"c2",X"ba",X"08",X"cd",X"fa",X"08", -- 0d60
  X"cd",X"23",X"0d",X"cd",X"7d",X"0d",X"f6",X"37", -- 0d68
  X"3a",X"f2",X"80",X"8f",X"b7",X"e8",X"c3",X"b0", -- 0d70
  X"04",X"cd",X"6c",X"07",X"28",X"2b",X"16",X"00", -- 0d78
  X"d5",X"0e",X"01",X"cd",X"7b",X"04",X"cd",X"f4", -- 0d80
  X"0d",X"22",X"15",X"81",X"2a",X"15",X"81",X"c1", -- 0d88
  X"78",X"fe",X"78",X"d4",X"6e",X"0d",X"7e",X"16", -- 0d90
  X"00",X"d6",X"b3",X"da",X"b5",X"0d",X"fe",X"03", -- 0d98
  X"d2",X"b5",X"0d",X"fe",X"01",X"17",X"aa",X"ba", -- 0da0
  X"57",X"da",X"9e",X"04",X"22",X"0a",X"81",X"cd", -- 0da8
  X"fa",X"08",X"c3",X"99",X"0d",X"7a",X"b7",X"c2", -- 0db0
  X"dd",X"0e",X"7e",X"22",X"0a",X"81",X"d6",X"ac", -- 0db8
  X"d8",X"fe",X"07",X"d0",X"5f",X"3a",X"f2",X"80", -- 0dc0
  X"3d",X"b3",X"7b",X"ca",X"3b",X"13",X"07",X"83", -- 0dc8
  X"5f",X"21",X"90",X"03",X"19",X"78",X"56",X"ba", -- 0dd0
  X"d0",X"23",X"cd",X"6e",X"0d",X"c5",X"01",X"8c", -- 0dd8
  X"0d",X"c5",X"43",X"4a",X"cd",X"81",X"17",X"58", -- 0de0
  X"51",X"4e",X"23",X"46",X"23",X"c5",X"2a",X"0a", -- 0de8
  X"81",X"c3",X"80",X"0d",X"af",X"32",X"f2",X"80", -- 0df0
  X"cd",X"fa",X"08",X"1e",X"24",X"ca",X"b2",X"04", -- 0df8
  X"da",X"57",X"18",X"cd",X"9c",X"09",X"d2",X"5c", -- 0e00
  X"0e",X"fe",X"26",X"c2",X"20",X"0e",X"cd",X"fa", -- 0e08
  X"08",X"fe",X"48",X"ca",X"a3",X"1c",X"fe",X"42", -- 0e10
  X"ca",X"1f",X"1d",X"1e",X"02",X"ca",X"b2",X"04", -- 0e18
  X"fe",X"ac",X"ca",X"f4",X"0d",X"fe",X"2e",X"ca", -- 0e20
  X"57",X"18",X"fe",X"ad",X"ca",X"4b",X"0e",X"fe", -- 0e28
  X"22",X"ca",X"04",X"12",X"fe",X"aa",X"ca",X"3d", -- 0e30
  X"0f",X"fe",X"a7",X"ca",X"68",X"11",X"d6",X"b6", -- 0e38
  X"d2",X"6d",X"0e",X"cd",X"79",X"0d",X"cd",X"6c", -- 0e40
  X"07",X"29",X"c9",X"16",X"7d",X"cd",X"80",X"0d", -- 0e48
  X"2a",X"15",X"81",X"e5",X"cd",X"79",X"17",X"cd", -- 0e50
  X"6e",X"0d",X"e1",X"c9",X"cd",X"62",X"0f",X"e5", -- 0e58
  X"eb",X"22",X"29",X"81",X"3a",X"f2",X"80",X"b7", -- 0e60
  X"cc",X"8e",X"17",X"e1",X"c9",X"06",X"00",X"07", -- 0e68
  X"4f",X"c5",X"cd",X"fa",X"08",X"79",X"fe",X"31", -- 0e70
  X"da",X"94",X"0e",X"cd",X"79",X"0d",X"cd",X"6c", -- 0e78
  X"07",X"2c",X"cd",X"6f",X"0d",X"eb",X"2a",X"29", -- 0e80
  X"81",X"e3",X"e5",X"eb",X"cd",X"cf",X"14",X"eb", -- 0e88
  X"e3",X"c3",X"9c",X"0e",X"cd",X"43",X"0e",X"e3", -- 0e90
  X"11",X"57",X"0e",X"d5",X"01",X"ef",X"01",X"09", -- 0e98
  X"4e",X"23",X"66",X"69",X"e9",X"15",X"fe",X"ad", -- 0ea0
  X"c8",X"fe",X"2d",X"c8",X"14",X"fe",X"2b",X"c8", -- 0ea8
  X"fe",X"ac",X"c8",X"2b",X"c9",X"f6",X"af",X"f5", -- 0eb0
  X"cd",X"6e",X"0d",X"cd",X"b0",X"09",X"f1",X"eb", -- 0eb8
  X"c1",X"e3",X"eb",X"cd",X"91",X"17",X"f5",X"cd", -- 0ec0
  X"b0",X"09",X"f1",X"c1",X"79",X"21",X"26",X"11", -- 0ec8
  X"c2",X"d8",X"0e",X"a3",X"4f",X"78",X"a2",X"e9", -- 0ed0
  X"b3",X"4f",X"78",X"b2",X"e9",X"21",X"ef",X"0e", -- 0ed8
  X"3a",X"f2",X"80",X"1f",X"7a",X"17",X"5f",X"16", -- 0ee0
  X"64",X"78",X"ba",X"d0",X"c3",X"dd",X"0d",X"f1", -- 0ee8
  X"0e",X"79",X"b7",X"1f",X"c1",X"d1",X"f5",X"cd", -- 0ef0
  X"70",X"0d",X"21",X"33",X"0f",X"e5",X"ca",X"cb", -- 0ef8
  X"17",X"af",X"32",X"f2",X"80",X"d5",X"cd",X"88", -- 0f00
  X"13",X"7e",X"23",X"23",X"4e",X"23",X"46",X"d1", -- 0f08
  X"c5",X"f5",X"cd",X"8c",X"13",X"cd",X"9f",X"17", -- 0f10
  X"f1",X"57",X"e1",X"7b",X"b2",X"c8",X"7a",X"d6", -- 0f18
  X"01",X"d8",X"af",X"bb",X"3c",X"d0",X"15",X"1d", -- 0f20
  X"0a",X"be",X"23",X"03",X"ca",X"1b",X"0f",X"3f", -- 0f28
  X"c3",X"5b",X"17",X"3c",X"8f",X"c1",X"a0",X"c6", -- 0f30
  X"ff",X"9f",X"c3",X"62",X"17",X"16",X"5a",X"cd", -- 0f38
  X"80",X"0d",X"cd",X"6e",X"0d",X"cd",X"b0",X"09", -- 0f40
  X"7b",X"2f",X"4f",X"7a",X"2f",X"cd",X"26",X"11", -- 0f48
  X"c1",X"c3",X"8c",X"0d",X"2b",X"cd",X"fa",X"08", -- 0f50
  X"c8",X"cd",X"6c",X"07",X"2c",X"01",X"54",X"0f", -- 0f58
  X"c5",X"f6",X"af",X"32",X"f1",X"80",X"46",X"cd", -- 0f60
  X"9c",X"09",X"da",X"9e",X"04",X"af",X"4f",X"32", -- 0f68
  X"f2",X"80",X"cd",X"fa",X"08",X"da",X"7e",X"0f", -- 0f70
  X"cd",X"9c",X"09",X"da",X"8b",X"0f",X"4f",X"cd", -- 0f78
  X"fa",X"08",X"da",X"7f",X"0f",X"cd",X"9c",X"09", -- 0f80
  X"d2",X"7f",X"0f",X"d6",X"24",X"c2",X"9a",X"0f", -- 0f88
  X"3c",X"32",X"f2",X"80",X"0f",X"81",X"4f",X"cd", -- 0f90
  X"fa",X"08",X"3a",X"10",X"81",X"3d",X"ca",X"47", -- 0f98
  X"10",X"f2",X"aa",X"0f",X"7e",X"d6",X"28",X"ca", -- 0fa0
  X"1f",X"10",X"af",X"32",X"10",X"81",X"e5",X"50", -- 0fa8
  X"59",X"2a",X"23",X"81",X"cd",X"66",X"07",X"11", -- 0fb0
  X"25",X"81",X"ca",X"91",X"16",X"2a",X"1d",X"81", -- 0fb8
  X"eb",X"2a",X"1b",X"81",X"cd",X"66",X"07",X"ca", -- 0fc0
  X"dd",X"0f",X"79",X"96",X"23",X"c2",X"d2",X"0f", -- 0fc8
  X"78",X"96",X"23",X"ca",X"11",X"10",X"23",X"23", -- 0fd0
  X"23",X"23",X"c3",X"c4",X"0f",X"e1",X"e3",X"d5", -- 0fd8
  X"11",X"5f",X"0e",X"cd",X"66",X"07",X"d1",X"ca", -- 0fe0
  X"14",X"10",X"e3",X"e5",X"c5",X"01",X"06",X"00", -- 0fe8
  X"2a",X"1f",X"81",X"e5",X"09",X"c1",X"e5",X"cd", -- 0ff0
  X"6a",X"04",X"e1",X"22",X"1f",X"81",X"60",X"69", -- 0ff8
  X"22",X"1d",X"81",X"2b",X"36",X"00",X"cd",X"66", -- 1000
  X"07",X"c2",X"03",X"10",X"d1",X"73",X"23",X"72", -- 1008
  X"23",X"eb",X"e1",X"c9",X"32",X"2c",X"81",X"21", -- 1010
  X"3a",X"04",X"22",X"29",X"81",X"e1",X"c9",X"e5", -- 1018
  X"2a",X"f1",X"80",X"e3",X"57",X"d5",X"c5",X"cd", -- 1020
  X"a4",X"09",X"c1",X"f1",X"eb",X"e3",X"e5",X"eb", -- 1028
  X"3c",X"57",X"7e",X"fe",X"2c",X"ca",X"25",X"10", -- 1030
  X"cd",X"6c",X"07",X"29",X"22",X"15",X"81",X"e1", -- 1038
  X"22",X"f1",X"80",X"1e",X"00",X"d5",X"11",X"e5", -- 1040
  X"f5",X"2a",X"1d",X"81",X"3e",X"19",X"eb",X"2a", -- 1048
  X"1f",X"81",X"eb",X"cd",X"66",X"07",X"ca",X"7f", -- 1050
  X"10",X"7e",X"b9",X"23",X"c2",X"61",X"10",X"7e", -- 1058
  X"b8",X"23",X"5e",X"23",X"56",X"23",X"c2",X"4d", -- 1060
  X"10",X"3a",X"f1",X"80",X"b7",X"c2",X"a7",X"04", -- 1068
  X"f1",X"44",X"4d",X"ca",X"91",X"16",X"96",X"ca", -- 1070
  X"dd",X"10",X"1e",X"10",X"c3",X"b2",X"04",X"11", -- 1078
  X"04",X"00",X"f1",X"ca",X"c5",X"09",X"71",X"23", -- 1080
  X"70",X"23",X"4f",X"cd",X"7b",X"04",X"23",X"23", -- 1088
  X"22",X"0a",X"81",X"71",X"23",X"3a",X"f1",X"80", -- 1090
  X"17",X"79",X"01",X"0b",X"00",X"d2",X"a2",X"10", -- 1098
  X"c1",X"03",X"71",X"23",X"70",X"23",X"f5",X"e5", -- 10a0
  X"cd",X"3c",X"18",X"eb",X"e1",X"f1",X"3d",X"c2", -- 10a8
  X"9a",X"10",X"f5",X"42",X"4b",X"eb",X"19",X"da", -- 10b0
  X"93",X"04",X"cd",X"84",X"04",X"22",X"1f",X"81", -- 10b8
  X"2b",X"36",X"00",X"cd",X"66",X"07",X"c2",X"c0", -- 10c0
  X"10",X"03",X"57",X"2a",X"0a",X"81",X"5e",X"eb", -- 10c8
  X"29",X"09",X"eb",X"2b",X"2b",X"73",X"23",X"72", -- 10d0
  X"23",X"f1",X"da",X"01",X"11",X"47",X"4f",X"7e", -- 10d8
  X"23",X"16",X"e1",X"5e",X"23",X"56",X"23",X"e3", -- 10e0
  X"f5",X"cd",X"66",X"07",X"d2",X"7a",X"10",X"e5", -- 10e8
  X"cd",X"3c",X"18",X"d1",X"19",X"f1",X"3d",X"44", -- 10f0
  X"4d",X"c2",X"e2",X"10",X"29",X"29",X"c1",X"09", -- 10f8
  X"eb",X"2a",X"15",X"81",X"c9",X"2a",X"1f",X"81", -- 1100
  X"eb",X"21",X"00",X"00",X"39",X"3a",X"f2",X"80", -- 1108
  X"b7",X"ca",X"21",X"11",X"cd",X"88",X"13",X"cd", -- 1110
  X"88",X"12",X"2a",X"9f",X"80",X"eb",X"2a",X"08", -- 1118
  X"81",X"7d",X"93",X"4f",X"7c",X"9a",X"41",X"50", -- 1120
  X"1e",X"00",X"21",X"f2",X"80",X"73",X"06",X"90", -- 1128
  X"c3",X"67",X"17",X"3a",X"f0",X"80",X"47",X"af", -- 1130
  X"c3",X"27",X"11",X"cd",X"be",X"11",X"cd",X"b0", -- 1138
  X"11",X"01",X"95",X"0a",X"c5",X"d5",X"cd",X"6c", -- 1140
  X"07",X"28",X"cd",X"62",X"0f",X"e5",X"eb",X"2b", -- 1148
  X"56",X"2b",X"5e",X"e1",X"cd",X"6e",X"0d",X"cd", -- 1150
  X"6c",X"07",X"29",X"cd",X"6c",X"07",X"b4",X"44", -- 1158
  X"4d",X"e3",X"71",X"23",X"70",X"c3",X"fd",X"11", -- 1160
  X"cd",X"be",X"11",X"d5",X"cd",X"43",X"0e",X"cd", -- 1168
  X"6e",X"0d",X"e3",X"5e",X"23",X"56",X"23",X"7a", -- 1170
  X"b3",X"ca",X"aa",X"04",X"7e",X"23",X"66",X"6f", -- 1178
  X"e5",X"2a",X"23",X"81",X"e3",X"22",X"23",X"81", -- 1180
  X"2a",X"27",X"81",X"e5",X"2a",X"25",X"81",X"e5", -- 1188
  X"21",X"25",X"81",X"d5",X"cd",X"a8",X"17",X"e1", -- 1190
  X"cd",X"6b",X"0d",X"2b",X"cd",X"fa",X"08",X"c2", -- 1198
  X"9e",X"04",X"e1",X"22",X"25",X"81",X"e1",X"22", -- 11a0
  X"27",X"81",X"e1",X"22",X"23",X"81",X"e1",X"c9", -- 11a8
  X"e5",X"2a",X"a1",X"80",X"23",X"7c",X"b5",X"e1", -- 11b0
  X"c0",X"1e",X"16",X"c3",X"b2",X"04",X"cd",X"6c", -- 11b8
  X"07",X"a7",X"3e",X"80",X"32",X"10",X"81",X"b6", -- 11c0
  X"47",X"cd",X"67",X"0f",X"c3",X"6e",X"0d",X"cd", -- 11c8
  X"6e",X"0d",X"cd",X"f5",X"18",X"cd",X"03",X"12", -- 11d0
  X"cd",X"88",X"13",X"01",X"e3",X"13",X"c5",X"7e", -- 11d8
  X"23",X"23",X"e5",X"cd",X"5e",X"12",X"e1",X"4e", -- 11e0
  X"23",X"46",X"cd",X"f7",X"11",X"e5",X"6f",X"cd", -- 11e8
  X"7b",X"13",X"d1",X"c9",X"cd",X"5e",X"12",X"21", -- 11f0
  X"04",X"81",X"e5",X"77",X"23",X"23",X"73",X"23", -- 11f8
  X"72",X"e1",X"c9",X"2b",X"06",X"22",X"50",X"e5", -- 1200
  X"0e",X"ff",X"23",X"7e",X"0c",X"b7",X"ca",X"19", -- 1208
  X"12",X"ba",X"ca",X"19",X"12",X"b8",X"c2",X"0a", -- 1210
  X"12",X"fe",X"22",X"cc",X"fa",X"08",X"e3",X"23", -- 1218
  X"eb",X"79",X"cd",X"f7",X"11",X"11",X"04",X"81", -- 1220
  X"2a",X"f6",X"80",X"22",X"29",X"81",X"3e",X"01", -- 1228
  X"32",X"f2",X"80",X"cd",X"ab",X"17",X"cd",X"66", -- 1230
  X"07",X"22",X"f6",X"80",X"e1",X"7e",X"c0",X"1e", -- 1238
  X"1e",X"c3",X"b2",X"04",X"23",X"cd",X"03",X"12", -- 1240
  X"cd",X"88",X"13",X"cd",X"9f",X"17",X"1c",X"1d", -- 1248
  X"c8",X"0a",X"cd",X"77",X"07",X"fe",X"0d",X"cc", -- 1250
  X"b0",X"0b",X"03",X"c3",X"4f",X"12",X"b7",X"0e", -- 1258
  X"f1",X"f5",X"2a",X"9f",X"80",X"eb",X"2a",X"08", -- 1260
  X"81",X"2f",X"4f",X"06",X"ff",X"09",X"23",X"cd", -- 1268
  X"66",X"07",X"da",X"7c",X"12",X"22",X"08",X"81", -- 1270
  X"23",X"eb",X"f1",X"c9",X"f1",X"1e",X"1a",X"ca", -- 1278
  X"b2",X"04",X"bf",X"f5",X"01",X"60",X"12",X"c5", -- 1280
  X"2a",X"f4",X"80",X"22",X"08",X"81",X"21",X"00", -- 1288
  X"00",X"e5",X"2a",X"9f",X"80",X"e5",X"21",X"f8", -- 1290
  X"80",X"eb",X"2a",X"f6",X"80",X"eb",X"cd",X"66", -- 1298
  X"07",X"01",X"99",X"12",X"c2",X"ed",X"12",X"2a", -- 12a0
  X"1b",X"81",X"eb",X"2a",X"1d",X"81",X"eb",X"cd", -- 12a8
  X"66",X"07",X"ca",X"c0",X"12",X"7e",X"23",X"23", -- 12b0
  X"b7",X"cd",X"f0",X"12",X"c3",X"aa",X"12",X"c1", -- 12b8
  X"eb",X"2a",X"1f",X"81",X"eb",X"cd",X"66",X"07", -- 12c0
  X"ca",X"16",X"13",X"cd",X"9f",X"17",X"7b",X"e5", -- 12c8
  X"09",X"b7",X"f2",X"bf",X"12",X"22",X"0a",X"81", -- 12d0
  X"e1",X"4e",X"06",X"00",X"09",X"09",X"23",X"eb", -- 12d8
  X"2a",X"0a",X"81",X"eb",X"cd",X"66",X"07",X"ca", -- 12e0
  X"c0",X"12",X"01",X"df",X"12",X"c5",X"f6",X"80", -- 12e8
  X"7e",X"23",X"23",X"5e",X"23",X"56",X"23",X"f0", -- 12f0
  X"b7",X"c8",X"44",X"4d",X"2a",X"08",X"81",X"cd", -- 12f8
  X"66",X"07",X"60",X"69",X"d8",X"e1",X"e3",X"cd", -- 1300
  X"66",X"07",X"e3",X"e5",X"60",X"69",X"d0",X"c1", -- 1308
  X"f1",X"f1",X"e5",X"d5",X"c5",X"c9",X"d1",X"e1", -- 1310
  X"7d",X"b4",X"c8",X"2b",X"46",X"2b",X"4e",X"e5", -- 1318
  X"2b",X"2b",X"6e",X"26",X"00",X"09",X"50",X"59", -- 1320
  X"2b",X"44",X"4d",X"2a",X"08",X"81",X"cd",X"6d", -- 1328
  X"04",X"e1",X"71",X"23",X"70",X"69",X"60",X"2b", -- 1330
  X"c3",X"8b",X"12",X"c5",X"e5",X"2a",X"29",X"81", -- 1338
  X"e3",X"cd",X"f4",X"0d",X"e3",X"cd",X"6f",X"0d", -- 1340
  X"7e",X"e5",X"2a",X"29",X"81",X"e5",X"86",X"1e", -- 1348
  X"1c",X"da",X"b2",X"04",X"cd",X"f4",X"11",X"d1", -- 1350
  X"cd",X"8c",X"13",X"e3",X"cd",X"8b",X"13",X"e5", -- 1358
  X"2a",X"06",X"81",X"eb",X"cd",X"72",X"13",X"cd", -- 1360
  X"72",X"13",X"21",X"89",X"0d",X"e3",X"e5",X"c3", -- 1368
  X"25",X"12",X"e1",X"e3",X"7e",X"23",X"23",X"4e", -- 1370
  X"23",X"46",X"6f",X"2c",X"2d",X"c8",X"0a",X"12", -- 1378
  X"03",X"13",X"c3",X"7c",X"13",X"cd",X"6f",X"0d", -- 1380
  X"2a",X"29",X"81",X"eb",X"cd",X"a6",X"13",X"eb", -- 1388
  X"c0",X"d5",X"50",X"59",X"1b",X"4e",X"2a",X"08", -- 1390
  X"81",X"cd",X"66",X"07",X"c2",X"a4",X"13",X"47", -- 1398
  X"09",X"22",X"08",X"81",X"e1",X"c9",X"2a",X"f6", -- 13a0
  X"80",X"2b",X"46",X"2b",X"4e",X"2b",X"2b",X"cd", -- 13a8
  X"66",X"07",X"c0",X"22",X"f6",X"80",X"c9",X"01", -- 13b0
  X"36",X"11",X"c5",X"cd",X"85",X"13",X"af",X"57", -- 13b8
  X"32",X"f2",X"80",X"7e",X"b7",X"c9",X"01",X"36", -- 13c0
  X"11",X"c5",X"cd",X"bb",X"13",X"ca",X"c5",X"09", -- 13c8
  X"23",X"23",X"5e",X"23",X"56",X"1a",X"c9",X"3e", -- 13d0
  X"01",X"cd",X"f4",X"11",X"cd",X"d2",X"14",X"2a", -- 13d8
  X"06",X"81",X"73",X"c1",X"c3",X"25",X"12",X"cd", -- 13e0
  X"82",X"14",X"af",X"e3",X"4f",X"e5",X"7e",X"b8", -- 13e8
  X"da",X"f5",X"13",X"78",X"11",X"0e",X"00",X"c5", -- 13f0
  X"cd",X"5e",X"12",X"c1",X"e1",X"e5",X"23",X"23", -- 13f8
  X"46",X"23",X"66",X"68",X"06",X"00",X"09",X"44", -- 1400
  X"4d",X"cd",X"f7",X"11",X"6f",X"cd",X"7b",X"13", -- 1408
  X"d1",X"cd",X"8c",X"13",X"c3",X"25",X"12",X"cd", -- 1410
  X"82",X"14",X"d1",X"d5",X"1a",X"90",X"c3",X"eb", -- 1418
  X"13",X"eb",X"7e",X"cd",X"87",X"14",X"04",X"05", -- 1420
  X"ca",X"c5",X"09",X"c5",X"1e",X"ff",X"fe",X"29", -- 1428
  X"ca",X"3a",X"14",X"cd",X"6c",X"07",X"2c",X"cd", -- 1430
  X"cf",X"14",X"cd",X"6c",X"07",X"29",X"f1",X"e3", -- 1438
  X"01",X"ed",X"13",X"c5",X"3d",X"be",X"06",X"00", -- 1440
  X"d0",X"4f",X"7e",X"91",X"bb",X"47",X"d8",X"43", -- 1448
  X"c9",X"cd",X"bb",X"13",X"ca",X"70",X"15",X"5f", -- 1450
  X"23",X"23",X"7e",X"23",X"66",X"6f",X"e5",X"19", -- 1458
  X"46",X"72",X"e3",X"c5",X"7e",X"fe",X"24",X"c2", -- 1460
  X"70",X"14",X"cd",X"a3",X"1c",X"c3",X"7e",X"14", -- 1468
  X"fe",X"25",X"c2",X"7b",X"14",X"cd",X"1f",X"1d", -- 1470
  X"c3",X"7e",X"14",X"cd",X"57",X"18",X"c1",X"e1", -- 1478
  X"70",X"c9",X"eb",X"cd",X"6c",X"07",X"29",X"c1", -- 1480
  X"d1",X"c5",X"43",X"c9",X"cd",X"d2",X"14",X"32", -- 1488
  X"84",X"80",X"cd",X"83",X"80",X"c3",X"36",X"11", -- 1490
  X"cd",X"bc",X"14",X"c3",X"4b",X"80",X"cd",X"bc", -- 1498
  X"14",X"f5",X"1e",X"00",X"2b",X"cd",X"fa",X"08", -- 14a0
  X"ca",X"b2",X"14",X"cd",X"6c",X"07",X"2c",X"cd", -- 14a8
  X"cf",X"14",X"c1",X"cd",X"83",X"80",X"ab",X"a0", -- 14b0
  X"ca",X"b3",X"14",X"c9",X"cd",X"cf",X"14",X"32", -- 14b8
  X"84",X"80",X"32",X"4c",X"80",X"cd",X"6c",X"07", -- 14c0
  X"2c",X"c3",X"cf",X"14",X"cd",X"fa",X"08",X"cd", -- 14c8
  X"6b",X"0d",X"cd",X"aa",X"09",X"7a",X"b7",X"c2", -- 14d0
  X"c5",X"09",X"2b",X"cd",X"fa",X"08",X"7b",X"c9", -- 14d8
  X"cd",X"b0",X"09",X"1a",X"c3",X"36",X"11",X"cd", -- 14e0
  X"6b",X"0d",X"cd",X"b0",X"09",X"d5",X"cd",X"6c", -- 14e8
  X"07",X"2c",X"cd",X"cf",X"14",X"d1",X"12",X"c9", -- 14f0
  X"21",X"ce",X"19",X"cd",X"9f",X"17",X"c3",X"0a", -- 14f8
  X"15",X"cd",X"9f",X"17",X"21",X"c1",X"d1",X"cd", -- 1500
  X"79",X"17",X"78",X"b7",X"c8",X"3a",X"2c",X"81", -- 1508
  X"b7",X"ca",X"91",X"17",X"90",X"d2",X"24",X"15", -- 1510
  X"2f",X"3c",X"eb",X"cd",X"81",X"17",X"eb",X"cd", -- 1518
  X"91",X"17",X"c1",X"d1",X"fe",X"19",X"d0",X"f5", -- 1520
  X"cd",X"b6",X"17",X"67",X"f1",X"cd",X"cf",X"15", -- 1528
  X"b4",X"21",X"29",X"81",X"f2",X"4a",X"15",X"cd", -- 1530
  X"af",X"15",X"d2",X"90",X"15",X"23",X"34",X"ca", -- 1538
  X"ad",X"04",X"2e",X"01",X"cd",X"e5",X"15",X"c3", -- 1540
  X"90",X"15",X"af",X"90",X"47",X"7e",X"9b",X"5f", -- 1548
  X"23",X"7e",X"9a",X"57",X"23",X"7e",X"99",X"4f", -- 1550
  X"dc",X"bb",X"15",X"68",X"63",X"af",X"47",X"79", -- 1558
  X"b7",X"c2",X"7d",X"15",X"4a",X"54",X"65",X"6f", -- 1560
  X"78",X"d6",X"08",X"fe",X"e0",X"c2",X"5e",X"15", -- 1568
  X"af",X"32",X"2c",X"81",X"c9",X"05",X"29",X"7a", -- 1570
  X"17",X"57",X"79",X"8f",X"4f",X"f2",X"75",X"15", -- 1578
  X"78",X"5c",X"45",X"b7",X"ca",X"90",X"15",X"21", -- 1580
  X"2c",X"81",X"86",X"77",X"d2",X"70",X"15",X"c8", -- 1588
  X"78",X"21",X"2c",X"81",X"b7",X"fc",X"a2",X"15", -- 1590
  X"46",X"23",X"7e",X"e6",X"80",X"a9",X"4f",X"c3", -- 1598
  X"91",X"17",X"1c",X"c0",X"14",X"c0",X"0c",X"c0", -- 15a0
  X"0e",X"80",X"34",X"c0",X"c3",X"ad",X"04",X"7e", -- 15a8
  X"83",X"5f",X"23",X"7e",X"8a",X"57",X"23",X"7e", -- 15b0
  X"89",X"4f",X"c9",X"21",X"2d",X"81",X"7e",X"2f", -- 15b8
  X"77",X"af",X"6f",X"90",X"47",X"7d",X"9b",X"5f", -- 15c0
  X"7d",X"9a",X"57",X"7d",X"99",X"4f",X"c9",X"06", -- 15c8
  X"00",X"d6",X"08",X"da",X"de",X"15",X"43",X"5a", -- 15d0
  X"51",X"0e",X"00",X"c3",X"d1",X"15",X"c6",X"09", -- 15d8
  X"6f",X"af",X"2d",X"c8",X"79",X"1f",X"4f",X"7a", -- 15e0
  X"1f",X"57",X"7b",X"1f",X"5f",X"78",X"1f",X"47", -- 15e8
  X"c3",X"e1",X"15",X"00",X"00",X"00",X"81",X"03", -- 15f0
  X"aa",X"56",X"19",X"80",X"f1",X"22",X"76",X"80", -- 15f8
  X"45",X"aa",X"38",X"82",X"cd",X"50",X"17",X"b7", -- 1600
  X"ea",X"c5",X"09",X"21",X"2c",X"81",X"7e",X"01", -- 1608
  X"35",X"80",X"11",X"f3",X"04",X"90",X"f5",X"70", -- 1610
  X"d5",X"c5",X"cd",X"0a",X"15",X"c1",X"d1",X"04", -- 1618
  X"cd",X"a6",X"16",X"21",X"f3",X"15",X"cd",X"01", -- 1620
  X"15",X"21",X"f7",X"15",X"cd",X"98",X"1a",X"01", -- 1628
  X"80",X"80",X"11",X"00",X"00",X"cd",X"0a",X"15", -- 1630
  X"f1",X"cd",X"cb",X"18",X"01",X"31",X"80",X"11", -- 1638
  X"18",X"72",X"21",X"c1",X"d1",X"cd",X"50",X"17", -- 1640
  X"c8",X"2e",X"00",X"cd",X"0e",X"17",X"79",X"32", -- 1648
  X"3b",X"81",X"eb",X"22",X"3c",X"81",X"01",X"00", -- 1650
  X"00",X"50",X"58",X"21",X"5b",X"15",X"e5",X"21", -- 1658
  X"67",X"16",X"e5",X"e5",X"21",X"29",X"81",X"7e", -- 1660
  X"23",X"b7",X"ca",X"93",X"16",X"e5",X"2e",X"08", -- 1668
  X"1f",X"67",X"79",X"d2",X"81",X"16",X"e5",X"2a", -- 1670
  X"3c",X"81",X"19",X"eb",X"e1",X"3a",X"3b",X"81", -- 1678
  X"89",X"1f",X"4f",X"7a",X"1f",X"57",X"7b",X"1f", -- 1680
  X"5f",X"78",X"1f",X"47",X"2d",X"7c",X"c2",X"70", -- 1688
  X"16",X"e1",X"c9",X"43",X"5a",X"51",X"4f",X"c9", -- 1690
  X"cd",X"81",X"17",X"01",X"20",X"84",X"11",X"00", -- 1698
  X"00",X"cd",X"91",X"17",X"c1",X"d1",X"cd",X"50", -- 16a0
  X"17",X"ca",X"a1",X"04",X"2e",X"ff",X"cd",X"0e", -- 16a8
  X"17",X"34",X"34",X"2b",X"7e",X"32",X"57",X"80", -- 16b0
  X"2b",X"7e",X"32",X"53",X"80",X"2b",X"7e",X"32", -- 16b8
  X"4f",X"80",X"41",X"eb",X"af",X"4f",X"57",X"5f", -- 16c0
  X"32",X"5a",X"80",X"e5",X"c5",X"7d",X"cd",X"4e", -- 16c8
  X"80",X"de",X"00",X"3f",X"d2",X"de",X"16",X"32", -- 16d0
  X"5a",X"80",X"f1",X"f1",X"37",X"d2",X"c1",X"e1", -- 16d8
  X"79",X"3c",X"3d",X"1f",X"fa",X"91",X"15",X"17", -- 16e0
  X"7b",X"17",X"5f",X"7a",X"17",X"57",X"79",X"17", -- 16e8
  X"4f",X"29",X"78",X"17",X"47",X"3a",X"5a",X"80", -- 16f0
  X"17",X"32",X"5a",X"80",X"79",X"b2",X"b3",X"c2", -- 16f8
  X"cb",X"16",X"e5",X"21",X"2c",X"81",X"35",X"e1", -- 1700
  X"c2",X"cb",X"16",X"c3",X"ad",X"04",X"78",X"b7", -- 1708
  X"ca",X"32",X"17",X"7d",X"21",X"2c",X"81",X"ae", -- 1710
  X"80",X"47",X"1f",X"a8",X"78",X"f2",X"31",X"17", -- 1718
  X"c6",X"80",X"77",X"ca",X"91",X"16",X"cd",X"b6", -- 1720
  X"17",X"77",X"2b",X"c9",X"cd",X"50",X"17",X"2f", -- 1728
  X"e1",X"b7",X"e1",X"f2",X"70",X"15",X"c3",X"ad", -- 1730
  X"04",X"cd",X"9c",X"17",X"78",X"b7",X"c8",X"c6", -- 1738
  X"02",X"da",X"ad",X"04",X"47",X"cd",X"0a",X"15", -- 1740
  X"21",X"2c",X"81",X"34",X"c0",X"c3",X"ad",X"04", -- 1748
  X"3a",X"2c",X"81",X"b7",X"c8",X"3a",X"2b",X"81", -- 1750
  X"fe",X"2f",X"17",X"9f",X"c0",X"3c",X"c9",X"cd", -- 1758
  X"50",X"17",X"06",X"88",X"11",X"00",X"00",X"21", -- 1760
  X"2c",X"81",X"4f",X"70",X"06",X"00",X"23",X"36", -- 1768
  X"80",X"17",X"c3",X"58",X"15",X"cd",X"50",X"17", -- 1770
  X"f0",X"21",X"2b",X"81",X"7e",X"ee",X"80",X"77", -- 1778
  X"c9",X"eb",X"2a",X"29",X"81",X"e3",X"e5",X"2a", -- 1780
  X"2b",X"81",X"e3",X"e5",X"eb",X"c9",X"cd",X"9f", -- 1788
  X"17",X"eb",X"22",X"29",X"81",X"60",X"69",X"22", -- 1790
  X"2b",X"81",X"eb",X"c9",X"21",X"29",X"81",X"5e", -- 1798
  X"23",X"56",X"23",X"4e",X"23",X"46",X"23",X"c9", -- 17a0
  X"11",X"29",X"81",X"06",X"04",X"1a",X"77",X"13", -- 17a8
  X"23",X"05",X"c2",X"ad",X"17",X"c9",X"21",X"2b", -- 17b0
  X"81",X"7e",X"07",X"37",X"1f",X"77",X"3f",X"1f", -- 17b8
  X"23",X"23",X"77",X"79",X"07",X"37",X"1f",X"4f", -- 17c0
  X"1f",X"ae",X"c9",X"78",X"b7",X"ca",X"50",X"17", -- 17c8
  X"21",X"59",X"17",X"e5",X"cd",X"50",X"17",X"79", -- 17d0
  X"c8",X"21",X"2b",X"81",X"ae",X"79",X"f8",X"cd", -- 17d8
  X"e5",X"17",X"1f",X"a9",X"c9",X"23",X"78",X"be", -- 17e0
  X"c0",X"2b",X"79",X"be",X"c0",X"2b",X"7a",X"be", -- 17e8
  X"c0",X"2b",X"7b",X"96",X"c0",X"e1",X"e1",X"c9", -- 17f0
  X"47",X"4f",X"57",X"5f",X"b7",X"c8",X"e5",X"cd", -- 17f8
  X"9c",X"17",X"cd",X"b6",X"17",X"ae",X"67",X"fc", -- 1800
  X"1c",X"18",X"3e",X"98",X"90",X"cd",X"cf",X"15", -- 1808
  X"7c",X"17",X"dc",X"a2",X"15",X"06",X"00",X"dc", -- 1810
  X"bb",X"15",X"e1",X"c9",X"1b",X"7a",X"a3",X"3c", -- 1818
  X"c0",X"0b",X"c9",X"21",X"2c",X"81",X"7e",X"fe", -- 1820
  X"98",X"3a",X"29",X"81",X"d0",X"7e",X"cd",X"f8", -- 1828
  X"17",X"36",X"98",X"7b",X"f5",X"79",X"17",X"cd", -- 1830
  X"58",X"15",X"f1",X"c9",X"21",X"00",X"00",X"78", -- 1838
  X"b1",X"c8",X"3e",X"10",X"29",X"da",X"7a",X"10", -- 1840
  X"eb",X"29",X"eb",X"d2",X"52",X"18",X"09",X"da", -- 1848
  X"7a",X"10",X"3d",X"c2",X"44",X"18",X"c9",X"fe", -- 1850
  X"2d",X"f5",X"ca",X"63",X"18",X"fe",X"2b",X"ca", -- 1858
  X"63",X"18",X"2b",X"cd",X"70",X"15",X"47",X"57", -- 1860
  X"5f",X"2f",X"4f",X"cd",X"fa",X"08",X"da",X"b4", -- 1868
  X"18",X"fe",X"2e",X"ca",X"8f",X"18",X"fe",X"45", -- 1870
  X"c2",X"93",X"18",X"cd",X"fa",X"08",X"cd",X"a5", -- 1878
  X"0e",X"cd",X"fa",X"08",X"da",X"d6",X"18",X"14", -- 1880
  X"c2",X"93",X"18",X"af",X"93",X"5f",X"0c",X"0c", -- 1888
  X"ca",X"6b",X"18",X"e5",X"7b",X"90",X"f4",X"ac", -- 1890
  X"18",X"f2",X"a2",X"18",X"f5",X"cd",X"98",X"16", -- 1898
  X"f1",X"3c",X"c2",X"96",X"18",X"d1",X"f1",X"cc", -- 18a0
  X"79",X"17",X"eb",X"c9",X"c8",X"f5",X"cd",X"39", -- 18a8
  X"17",X"f1",X"3d",X"c9",X"d5",X"57",X"78",X"89", -- 18b0
  X"47",X"c5",X"e5",X"d5",X"cd",X"39",X"17",X"f1", -- 18b8
  X"d6",X"30",X"cd",X"cb",X"18",X"e1",X"c1",X"d1", -- 18c0
  X"c3",X"6b",X"18",X"cd",X"81",X"17",X"cd",X"62", -- 18c8
  X"17",X"c1",X"d1",X"c3",X"0a",X"15",X"7b",X"07", -- 18d0
  X"07",X"83",X"07",X"86",X"d6",X"30",X"5f",X"c3", -- 18d8
  X"81",X"18",X"e5",X"21",X"36",X"04",X"cd",X"45", -- 18e0
  X"12",X"e1",X"eb",X"af",X"06",X"98",X"cd",X"67", -- 18e8
  X"17",X"21",X"44",X"12",X"e5",X"21",X"2e",X"81", -- 18f0
  X"e5",X"cd",X"50",X"17",X"36",X"20",X"f2",X"03", -- 18f8
  X"19",X"36",X"2d",X"23",X"36",X"30",X"ca",X"b9", -- 1900
  X"19",X"e5",X"fc",X"79",X"17",X"af",X"f5",X"cd", -- 1908
  X"bf",X"19",X"01",X"43",X"91",X"11",X"f8",X"4f", -- 1910
  X"cd",X"cb",X"17",X"b7",X"e2",X"30",X"19",X"f1", -- 1918
  X"cd",X"ad",X"18",X"f5",X"c3",X"12",X"19",X"cd", -- 1920
  X"98",X"16",X"f1",X"3c",X"f5",X"cd",X"bf",X"19", -- 1928
  X"cd",X"f8",X"14",X"3c",X"cd",X"f8",X"17",X"cd", -- 1930
  X"91",X"17",X"01",X"06",X"03",X"f1",X"81",X"3c", -- 1938
  X"fa",X"4c",X"19",X"fe",X"08",X"d2",X"4c",X"19", -- 1940
  X"3c",X"47",X"3e",X"02",X"3d",X"3d",X"e1",X"f5", -- 1948
  X"11",X"d2",X"19",X"05",X"c2",X"5d",X"19",X"36", -- 1950
  X"2e",X"23",X"36",X"30",X"23",X"05",X"36",X"2e", -- 1958
  X"cc",X"a6",X"17",X"c5",X"e5",X"d5",X"cd",X"9c", -- 1960
  X"17",X"e1",X"06",X"2f",X"04",X"7b",X"96",X"5f", -- 1968
  X"23",X"7a",X"9e",X"57",X"23",X"79",X"9e",X"4f", -- 1970
  X"2b",X"2b",X"d2",X"6c",X"19",X"cd",X"af",X"15", -- 1978
  X"23",X"cd",X"91",X"17",X"eb",X"e1",X"70",X"23", -- 1980
  X"c1",X"0d",X"c2",X"5d",X"19",X"05",X"ca",X"9d", -- 1988
  X"19",X"2b",X"7e",X"fe",X"30",X"ca",X"91",X"19", -- 1990
  X"fe",X"2e",X"c4",X"a6",X"17",X"f1",X"ca",X"bc", -- 1998
  X"19",X"36",X"45",X"23",X"36",X"2b",X"f2",X"ad", -- 19a0
  X"19",X"36",X"2d",X"2f",X"3c",X"06",X"2f",X"04", -- 19a8
  X"d6",X"0a",X"d2",X"af",X"19",X"c6",X"3a",X"23", -- 19b0
  X"70",X"23",X"77",X"23",X"71",X"e1",X"c9",X"01", -- 19b8
  X"74",X"94",X"11",X"f7",X"23",X"cd",X"cb",X"17", -- 19c0
  X"b7",X"e1",X"e2",X"27",X"19",X"e9",X"00",X"00", -- 19c8
  X"00",X"80",X"a0",X"86",X"01",X"10",X"27",X"00", -- 19d0
  X"e8",X"03",X"00",X"64",X"00",X"00",X"0a",X"00", -- 19d8
  X"00",X"01",X"00",X"00",X"21",X"79",X"17",X"e3", -- 19e0
  X"e9",X"cd",X"81",X"17",X"21",X"ce",X"19",X"cd", -- 19e8
  X"8e",X"17",X"c1",X"d1",X"cd",X"50",X"17",X"78", -- 19f0
  X"ca",X"37",X"1a",X"f2",X"02",X"1a",X"b7",X"ca", -- 19f8
  X"a1",X"04",X"b7",X"ca",X"71",X"15",X"d5",X"c5", -- 1a00
  X"79",X"f6",X"7f",X"cd",X"9c",X"17",X"f2",X"1f", -- 1a08
  X"1a",X"d5",X"c5",X"cd",X"23",X"18",X"c1",X"d1", -- 1a10
  X"f5",X"cd",X"cb",X"17",X"e1",X"7c",X"1f",X"e1", -- 1a18
  X"22",X"2b",X"81",X"e1",X"22",X"29",X"81",X"dc", -- 1a20
  X"e4",X"19",X"cc",X"79",X"17",X"d5",X"c5",X"cd", -- 1a28
  X"04",X"16",X"c1",X"d1",X"cd",X"45",X"16",X"cd", -- 1a30
  X"81",X"17",X"01",X"38",X"81",X"11",X"3b",X"aa", -- 1a38
  X"cd",X"45",X"16",X"3a",X"2c",X"81",X"fe",X"88", -- 1a40
  X"d2",X"2c",X"17",X"cd",X"23",X"18",X"c6",X"80", -- 1a48
  X"c6",X"02",X"da",X"2c",X"17",X"f5",X"21",X"f3", -- 1a50
  X"15",X"cd",X"fb",X"14",X"cd",X"3c",X"16",X"f1", -- 1a58
  X"c1",X"d1",X"f5",X"cd",X"07",X"15",X"cd",X"79", -- 1a60
  X"17",X"21",X"77",X"1a",X"cd",X"a7",X"1a",X"11", -- 1a68
  X"00",X"00",X"c1",X"4a",X"c3",X"45",X"16",X"08", -- 1a70
  X"40",X"2e",X"94",X"74",X"70",X"4f",X"2e",X"77", -- 1a78
  X"6e",X"02",X"88",X"7a",X"e6",X"a0",X"2a",X"7c", -- 1a80
  X"50",X"aa",X"aa",X"7e",X"ff",X"ff",X"7f",X"7f", -- 1a88
  X"00",X"00",X"80",X"81",X"00",X"00",X"00",X"81", -- 1a90
  X"cd",X"81",X"17",X"11",X"43",X"16",X"d5",X"e5", -- 1a98
  X"cd",X"9c",X"17",X"cd",X"45",X"16",X"e1",X"cd", -- 1aa0
  X"81",X"17",X"7e",X"23",X"cd",X"8e",X"17",X"06", -- 1aa8
  X"f1",X"c1",X"d1",X"3d",X"c8",X"d5",X"c5",X"f5", -- 1ab0
  X"e5",X"cd",X"45",X"16",X"e1",X"cd",X"9f",X"17", -- 1ab8
  X"e5",X"cd",X"0a",X"15",X"e1",X"c3",X"b0",X"1a", -- 1ac0
  X"cd",X"50",X"17",X"21",X"5e",X"80",X"fa",X"29", -- 1ac8
  X"1b",X"21",X"7f",X"80",X"cd",X"8e",X"17",X"21", -- 1ad0
  X"5e",X"80",X"c8",X"86",X"e6",X"07",X"06",X"00", -- 1ad8
  X"77",X"23",X"87",X"87",X"4f",X"09",X"cd",X"9f", -- 1ae0
  X"17",X"cd",X"45",X"16",X"3a",X"5d",X"80",X"3c", -- 1ae8
  X"e6",X"03",X"06",X"00",X"fe",X"01",X"88",X"32", -- 1af0
  X"5d",X"80",X"21",X"2d",X"1b",X"87",X"87",X"4f", -- 1af8
  X"09",X"cd",X"fb",X"14",X"cd",X"9c",X"17",X"7b", -- 1b00
  X"59",X"ee",X"4f",X"4f",X"36",X"80",X"2b",X"46", -- 1b08
  X"36",X"80",X"21",X"5c",X"80",X"34",X"7e",X"d6", -- 1b10
  X"ab",X"c2",X"20",X"1b",X"77",X"0c",X"15",X"1c", -- 1b18
  X"cd",X"5b",X"15",X"21",X"7f",X"80",X"c3",X"a8", -- 1b20
  X"17",X"77",X"2b",X"77",X"2b",X"77",X"c3",X"04", -- 1b28
  X"1b",X"68",X"b1",X"46",X"68",X"99",X"e9",X"92", -- 1b30
  X"69",X"10",X"d1",X"75",X"68",X"21",X"87",X"1b", -- 1b38
  X"cd",X"fb",X"14",X"cd",X"81",X"17",X"01",X"49", -- 1b40
  X"83",X"11",X"db",X"0f",X"cd",X"91",X"17",X"c1", -- 1b48
  X"d1",X"cd",X"a6",X"16",X"cd",X"81",X"17",X"cd", -- 1b50
  X"23",X"18",X"c1",X"d1",X"cd",X"07",X"15",X"21", -- 1b58
  X"8b",X"1b",X"cd",X"01",X"15",X"cd",X"50",X"17", -- 1b60
  X"37",X"f2",X"73",X"1b",X"cd",X"f8",X"14",X"cd", -- 1b68
  X"50",X"17",X"b7",X"f5",X"f4",X"79",X"17",X"21", -- 1b70
  X"8b",X"1b",X"cd",X"fb",X"14",X"f1",X"d4",X"79", -- 1b78
  X"17",X"21",X"8f",X"1b",X"c3",X"98",X"1a",X"db", -- 1b80
  X"0f",X"49",X"81",X"00",X"00",X"00",X"7f",X"05", -- 1b88
  X"ba",X"d7",X"1e",X"86",X"64",X"26",X"99",X"87", -- 1b90
  X"58",X"34",X"23",X"87",X"e0",X"5d",X"a5",X"86", -- 1b98
  X"da",X"0f",X"49",X"83",X"cd",X"81",X"17",X"cd", -- 1ba0
  X"43",X"1b",X"c1",X"e1",X"cd",X"81",X"17",X"eb", -- 1ba8
  X"cd",X"91",X"17",X"cd",X"3d",X"1b",X"c3",X"a4", -- 1bb0
  X"16",X"cd",X"50",X"17",X"fc",X"e4",X"19",X"fc", -- 1bb8
  X"79",X"17",X"3a",X"2c",X"81",X"fe",X"81",X"da", -- 1bc0
  X"d6",X"1b",X"01",X"00",X"81",X"51",X"59",X"cd", -- 1bc8
  X"a6",X"16",X"21",X"01",X"15",X"e5",X"21",X"e0", -- 1bd0
  X"1b",X"cd",X"98",X"1a",X"21",X"87",X"1b",X"c9", -- 1bd8
  X"09",X"4a",X"d7",X"3b",X"78",X"02",X"6e",X"84", -- 1be0
  X"7b",X"fe",X"c1",X"2f",X"7c",X"74",X"31",X"9a", -- 1be8
  X"7d",X"84",X"3d",X"5a",X"7d",X"c8",X"7f",X"91", -- 1bf0
  X"7e",X"e4",X"bb",X"4c",X"7e",X"6c",X"aa",X"aa", -- 1bf8
  X"7f",X"00",X"00",X"00",X"81",X"c9",X"d7",X"c9", -- 1c00
  X"3e",X"0c",X"c3",X"53",X"1d",X"cd",X"cf",X"14", -- 1c08
  X"7b",X"32",X"87",X"80",X"c9",X"cd",X"6b",X"0d", -- 1c10
  X"cd",X"b0",X"09",X"e5",X"d5",X"e1",X"22",X"8b", -- 1c18
  X"80",X"22",X"8d",X"80",X"e1",X"c9",X"cd",X"b0", -- 1c20
  X"09",X"d5",X"e1",X"46",X"23",X"7e",X"c3",X"27", -- 1c28
  X"11",X"cd",X"6b",X"0d",X"cd",X"b0",X"09",X"d5", -- 1c30
  X"cd",X"6c",X"07",X"2c",X"cd",X"6b",X"0d",X"cd", -- 1c38
  X"b0",X"09",X"e3",X"73",X"23",X"72",X"e1",X"c9", -- 1c40
  X"cd",X"6e",X"0d",X"cd",X"b0",X"09",X"c5",X"21", -- 1c48
  X"2e",X"81",X"7a",X"fe",X"00",X"ca",X"65",X"1c", -- 1c50
  X"cd",X"84",X"1c",X"78",X"fe",X"30",X"ca",X"63", -- 1c58
  X"1c",X"70",X"23",X"71",X"23",X"7b",X"cd",X"84", -- 1c60
  X"1c",X"7a",X"fe",X"00",X"c2",X"75",X"1c",X"78", -- 1c68
  X"fe",X"30",X"ca",X"77",X"1c",X"70",X"23",X"71", -- 1c70
  X"23",X"af",X"77",X"23",X"77",X"c1",X"21",X"2e", -- 1c78
  X"81",X"c3",X"d5",X"11",X"47",X"e6",X"0f",X"fe", -- 1c80
  X"0a",X"da",X"8e",X"1c",X"c6",X"07",X"c6",X"30", -- 1c88
  X"4f",X"78",X"0f",X"0f",X"0f",X"0f",X"e6",X"0f", -- 1c90
  X"fe",X"0a",X"da",X"9f",X"1c",X"c6",X"07",X"c6", -- 1c98
  X"30",X"47",X"c9",X"eb",X"21",X"00",X"00",X"cd", -- 1ca0
  X"bf",X"1c",X"da",X"e0",X"1c",X"c3",X"b6",X"1c", -- 1ca8
  X"cd",X"bf",X"1c",X"da",X"d7",X"1c",X"29",X"29", -- 1cb0
  X"29",X"29",X"b5",X"6f",X"c3",X"b0",X"1c",X"13", -- 1cb8
  X"1a",X"fe",X"20",X"ca",X"bf",X"1c",X"d6",X"30", -- 1cc0
  X"d8",X"fe",X"0a",X"da",X"d3",X"1c",X"d6",X"07", -- 1cc8
  X"fe",X"0a",X"d8",X"fe",X"10",X"3f",X"c9",X"eb", -- 1cd0
  X"7a",X"4b",X"e5",X"cd",X"26",X"11",X"e1",X"c9", -- 1cd8
  X"1e",X"26",X"c3",X"b2",X"04",X"cd",X"6e",X"0d", -- 1ce0
  X"cd",X"b0",X"09",X"c5",X"21",X"2e",X"81",X"06", -- 1ce8
  X"11",X"05",X"78",X"fe",X"01",X"ca",X"04",X"1d", -- 1cf0
  X"7b",X"17",X"5f",X"7a",X"17",X"57",X"d2",X"f1", -- 1cf8
  X"1c",X"c3",X"0a",X"1d",X"7b",X"17",X"5f",X"7a", -- 1d00
  X"17",X"57",X"3e",X"30",X"ce",X"00",X"77",X"23", -- 1d08
  X"05",X"c2",X"04",X"1d",X"af",X"77",X"23",X"77", -- 1d10
  X"c1",X"21",X"2e",X"81",X"c3",X"d5",X"11",X"eb", -- 1d18
  X"21",X"00",X"00",X"cd",X"3d",X"1d",X"da",X"4b", -- 1d20
  X"1d",X"d6",X"30",X"29",X"b5",X"6f",X"cd",X"3d", -- 1d28
  X"1d",X"d2",X"29",X"1d",X"eb",X"7a",X"4b",X"e5", -- 1d30
  X"cd",X"26",X"11",X"e1",X"c9",X"13",X"1a",X"fe", -- 1d38
  X"20",X"ca",X"3d",X"1d",X"fe",X"30",X"d8",X"fe", -- 1d40
  X"32",X"3f",X"c9",X"1e",X"28",X"c3",X"b2",X"04", -- 1d48
  X"c3",X"f1",X"00",X"c3",X"08",X"00",X"c3",X"00", -- 1d50
  X"00",X"3e",X"00",X"32",X"92",X"80",X"c3",X"f8", -- 1d58
  X"00",X"f5",X"a0",X"c1",X"b8",X"3e",X"00",X"c9", -- 1d60
  X"cd",X"77",X"07",X"c3",X"a6",X"0b",X"00",X"00", -- 1d68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1d98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1da0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1da8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1db0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1db8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1dc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1dc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1dd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1dd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1de0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1de8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1df0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1df8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1e98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ea0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ea8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1eb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1eb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ec0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ec8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ed0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ed8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ee0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ee8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ef0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ef8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1f98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fe0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1fe8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ff0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1ff8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2000
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2008
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2010
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2018
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2020
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2028
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2030
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2038
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2040
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2048
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2050
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2058
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2060
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2068
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2070
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2078
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2080
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2088
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2090
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2098
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 20f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2100
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2108
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2110
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2118
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2120
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2128
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2130
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2138
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2140
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2148
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2150
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2158
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2160
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2168
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2170
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2178
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2180
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2188
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2190
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2198
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 21f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2200
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2208
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2210
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2218
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2220
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2228
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2230
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2238
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2240
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2248
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2250
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2258
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2260
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2268
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2270
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2278
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2280
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2288
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2290
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2298
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 22f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2300
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2308
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2310
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2318
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2320
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2328
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2330
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2338
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2340
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2348
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2350
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2358
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2360
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2368
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2370
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2378
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2380
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2388
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2390
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2398
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 23f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2400
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2408
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2410
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2418
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2420
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2428
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2430
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2438
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2440
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2448
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2450
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2458
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2460
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2468
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2470
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2478
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2480
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2488
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2490
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2498
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 24f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2500
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2508
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2510
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2518
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2520
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2528
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2530
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2538
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2540
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2548
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2550
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2558
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2560
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2568
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2570
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2578
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2580
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2588
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2590
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2598
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 25f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2600
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2608
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2610
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2618
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2620
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2628
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2630
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2638
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2640
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2648
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2650
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2658
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2660
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2668
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2670
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2678
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2680
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2688
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2690
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2698
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 26f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2700
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2708
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2710
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2718
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2720
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2728
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2730
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2738
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2740
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2748
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2750
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2758
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2760
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2768
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2770
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2778
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2780
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2788
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2790
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2798
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 27f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2800
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2808
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2810
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2818
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2820
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2828
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2830
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2838
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2840
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2848
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2850
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2858
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2860
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2868
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2870
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2878
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2880
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2888
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2890
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2898
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 28f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2900
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2908
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2910
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2918
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2920
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2928
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2930
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2938
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2940
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2948
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2950
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2958
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2960
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2968
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2970
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2978
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2980
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2988
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2990
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2998
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 29f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2a98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2aa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2aa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ab0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ab8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ac0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ac8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ad0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ad8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ae0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ae8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2af0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2af8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2b98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ba0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ba8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2be0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2be8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2bf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2c98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ca0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ca8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ce0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ce8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2cf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2d98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2da0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2da8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2db0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2db8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2dd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2de0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2de8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2df0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2df8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2e98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ea0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ea8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2eb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2eb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ec0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ec8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ed0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ed8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ee0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ee8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ef0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ef8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2f98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fe0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2fe8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ff0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2ff8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3000
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3008
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3010
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3018
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3020
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3028
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3030
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3038
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3040
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3048
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3050
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3058
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3060
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3068
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3070
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3078
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3080
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3088
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3090
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3098
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 30f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3100
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3108
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3110
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3118
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3120
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3128
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3130
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3138
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3140
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3148
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3150
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3158
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3160
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3168
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3170
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3178
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3180
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3188
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3190
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3198
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 31f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3200
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3208
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3210
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3218
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3220
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3228
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3230
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3238
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3240
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3248
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3250
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3258
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3260
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3268
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3270
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3278
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3280
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3288
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3290
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3298
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 32f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3300
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3308
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3310
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3318
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3320
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3328
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3330
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3338
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3340
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3348
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3350
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3358
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3360
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3368
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3370
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3378
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3380
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3388
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3390
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3398
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 33f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3400
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3408
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3410
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3418
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3420
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3428
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3430
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3438
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3440
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3448
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3450
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3458
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3460
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3468
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3470
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3478
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3480
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3488
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3490
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3498
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 34f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3500
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3508
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3510
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3518
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3520
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3528
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3530
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3538
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3540
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3548
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3550
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3558
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3560
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3568
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3570
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3578
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3580
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3588
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3590
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3598
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 35f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3600
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3608
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3610
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3618
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3620
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3628
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3630
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3638
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3640
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3648
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3650
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3658
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3660
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3668
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3670
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3678
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3680
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3688
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3690
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3698
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 36f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3700
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3708
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3710
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3718
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3720
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3728
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3730
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3738
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3740
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3748
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3750
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3758
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3760
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3768
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3770
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3778
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3780
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3788
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3790
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3798
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 37f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3800
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3808
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3810
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3818
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3820
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3828
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3830
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3838
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3840
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3848
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3850
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3858
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3860
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3868
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3870
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3878
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3880
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3888
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3890
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3898
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 38f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3900
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3908
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3910
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3918
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3920
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3928
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3930
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3938
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3940
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3948
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3950
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3958
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3960
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3968
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3970
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3978
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3980
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3988
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3990
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3998
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39a0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39a8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39b0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39b8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39c0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39c8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39d0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39d8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39e0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39e8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39f0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 39f8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3a98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3aa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3aa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ab0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ab8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ac0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ac8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ad0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ad8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ae0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ae8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3af0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3af8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3b98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ba0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ba8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3be0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3be8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3bf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3c98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ca0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ca8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ce0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ce8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cf0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3cf8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3d98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3da0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3da8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3db0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3db8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3dd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3de0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3de8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3df0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3df8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3e98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ea0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ea8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3eb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3eb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ec0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ec8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ed0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ed8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ee0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ee8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ef0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ef8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f00
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f08
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f10
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f18
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f20
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f28
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f30
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f38
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f40
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f48
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f50
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f58
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f60
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f68
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f70
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f78
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f80
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f88
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f90
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3f98
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fa0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fa8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fb0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fb8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fc0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fc8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fd0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fd8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fe0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3fe8
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3ff0
  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"  -- 3ff8
  );

end package obj_code_pkg;
